module c880g( L1gat, L8gat, L13gat, L17gat, L26gat, L29gat, L36gat, L42gat, 
		L51gat, L55gat, L59gat, L68gat, L72gat, L73gat, L74gat, 
		L75gat, L80gat, L85gat, L86gat, L87gat, L88gat, L89gat, 
		L90gat, L91gat, L96gat, L101gat, L106gat, L111gat, L116gat, 
		L121gat, L126gat, L130gat, L135gat, L138gat, L143gat, L146gat, 
		L149gat, L152gat, L153gat, L156gat, L159gat, L165gat, L171gat, 
		L177gat, L183gat, L189gat, L195gat, L201gat, L207gat, L210gat, 
		L219gat, L228gat, L237gat, L246gat, L255gat, L259gat, L260gat, 
		L261gat, L267gat, L268gat, 
		L388gat, L389gat, L390gat, L391gat, L418gat, L419gat, L420gat, L421gat, 
		L422gat, L423gat, L446gat, L447gat, L448gat, L449gat, L450gat, 
		L767gat, L768gat, L850gat, L863gat, L864gat, L865gat, L866gat, 
		L874gat, L878gat, L879gat, L880gat );
input L1gat, L8gat, L13gat, L17gat, L26gat, L29gat, L36gat, L42gat, 
	L51gat, L55gat, L59gat, L68gat, L72gat, L73gat, L74gat, 
	L75gat, L80gat, L85gat, L86gat, L87gat, L88gat, L89gat, 
	L90gat, L91gat, L96gat, L101gat, L106gat, L111gat, L116gat, 
	L121gat, L126gat, L130gat, L135gat, L138gat, L143gat, L146gat, 
	L149gat, L152gat, L153gat, L156gat, L159gat, L165gat, L171gat, 
	L177gat, L183gat, L189gat, L195gat, L201gat, L207gat, L210gat, 
	L219gat, L228gat, L237gat, L246gat, L255gat, L259gat, L260gat, 
	L261gat, L267gat, L268gat ;
output L388gat, L389gat, L390gat, L391gat, L418gat, L419gat, L420gat, L421gat, 
	L422gat, L423gat, L446gat, L447gat, L448gat, L449gat, L450gat, 
	L767gat, L768gat, L850gat, L863gat, L864gat, L865gat, L866gat, 
	L874gat, L878gat, L879gat, L880gat ;




   NA4 U1 ( L1gat, L8gat, L13gat, L17gat, L269gat ); 
   NA4 U2 ( L1gat, L26gat, L13gat, L17gat, L270gat ); 
   AND3 U3 ( L29gat, L36gat, L42gat, L273gat ); 
   AND3 U4 ( L1gat, L26gat, L51gat, L276gat ); 
   NA4 U5 ( L1gat, L8gat, L51gat, L17gat, L279gat ); 
   NA4 U6 ( L1gat, L8gat, L13gat, L55gat, L280gat ); 
   NA4 U7 ( L59gat, L42gat, L68gat, L72gat, L284gat ); 
   NA2 U8 ( L29gat, L68gat, L285gat ); 
   NA3 U9 ( L59gat, L68gat, L74gat, L286gat ); 
   AND3 U10 ( L29gat, L75gat, L80gat, L287gat ); 
   AND3 U11 ( L29gat, L75gat, L42gat, L290gat ); 
   AND3 U12 ( L29gat, L36gat, L80gat, L291gat ); 
   AND3 U13 ( L29gat, L36gat, L42gat, L292gat ); 
   AND3 U14 ( L59gat, L75gat, L80gat, L293gat ); 
   AND3 U15 ( L59gat, L75gat, L42gat, L294gat ); 
   AND3 U16 ( L59gat, L36gat, L80gat, L295gat ); 
   AND3 U17 ( L59gat, L36gat, L42gat, L296gat ); 
   AND2 U18 ( L85gat, L86gat, L297gat ); 
   OR2 U19 ( L87gat, L88gat, L298gat ); 
   NA2 U20 ( L91gat, L96gat, L301gat ); 
   OR2 U21 ( L91gat, L96gat, L302gat ); 
   NA2 U22 ( L101gat, L106gat, L303gat ); 
   OR2 U23 ( L101gat, L106gat, L304gat ); 
   NA2 U24 ( L111gat, L116gat, L305gat ); 
   OR2 U25 ( L111gat, L116gat, L306gat ); 
   NA2 U26 ( L121gat, L126gat, L307gat ); 
   OR2 U27 ( L121gat, L126gat, L308gat ); 
   AND2 U28 ( L8gat, L138gat, L309gat ); 
   IN1 U29 ( L268gat, L310gat ); 
   AND2 U30 ( L51gat, L138gat, L316gat ); 
   AND2 U31 ( L17gat, L138gat, L317gat ); 
   AND2 U32 ( L152gat, L138gat, L318gat ); 
   NA2 U33 ( L59gat, L156gat, L319gat ); 
   NO2 U34 ( L17gat, L42gat, L322gat ); 
   AND2 U35 ( L17gat, L42gat, L323gat ); 
   NA2 U36 ( L159gat, L165gat, L324gat ); 
   OR2 U37 ( L159gat, L165gat, L325gat ); 
   NA2 U38 ( L171gat, L177gat, L326gat ); 
   OR2 U39 ( L171gat, L177gat, L327gat ); 
   NA2 U40 ( L183gat, L189gat, L328gat ); 
   OR2 U41 ( L183gat, L189gat, L329gat ); 
   NA2 U42 ( L195gat, L201gat, L330gat ); 
   OR2 U43 ( L195gat, L201gat, L331gat ); 
   AND2 U44 ( L210gat, L91gat, L332gat ); 
   AND2 U45 ( L210gat, L96gat, L333gat ); 
   AND2 U46 ( L210gat, L101gat, L334gat ); 
   AND2 U47 ( L210gat, L106gat, L335gat ); 
   AND2 U48 ( L210gat, L111gat, L336gat ); 
   AND2 U49 ( L255gat, L259gat, L337gat ); 
   AND2 U50 ( L210gat, L116gat, L338gat ); 
   AND2 U51 ( L255gat, L260gat, L339gat ); 
   AND2 U52 ( L210gat, L121gat, L340gat ); 
   AND2 U53 ( L255gat, L267gat, L341gat ); 
   IN1 U54 ( L269gat, L342gat ); 
   IN1 U55 ( L273gat, L343gat ); 
   OR2 U56 ( L270gat, L273gat, L344gat ); 
   IN1 U57 ( L276gat, L345gat ); 
   IN1 U58 ( L276gat, L346gat ); 
   IN1 U59 ( L279gat, L347gat ); 
   NO2 U60 ( L280gat, L284gat, L348gat ); 
   OR2 U61 ( L280gat, L285gat, L349gat ); 
   OR2 U62 ( L280gat, L286gat, L350gat ); 
   IN1 U63 ( L293gat, L351gat ); 
   IN1 U64 ( L294gat, L352gat ); 
   IN1 U65 ( L295gat, L353gat ); 
   IN1 U66 ( L296gat, L354gat ); 
   NA2 U67 ( L89gat, L298gat, L355gat ); 
   AND2 U68 ( L90gat, L298gat, L356gat ); 
   NA2 U69 ( L301gat, L302gat, L357gat ); 
   NA2 U70 ( L303gat, L304gat, L360gat ); 
   NA2 U71 ( L305gat, L306gat, L363gat ); 
   NA2 U72 ( L307gat, L308gat, L366gat ); 
   IN1 U73 ( L310gat, L369gat ); 
   NO2 U74 ( L322gat, L323gat, L375gat ); 
   NA2 U75 ( L324gat, L325gat, L376gat ); 
   NA2 U76 ( L326gat, L327gat, L379gat ); 
   NA2 U77 ( L328gat, L329gat, L382gat ); 
   NA2 U78 ( L330gat, L331gat, L385gat ); 
   BU1 U79 ( L290gat, L388gat ); 
   BU1 U80 ( L291gat, L389gat ); 
   BU1 U81 ( L292gat, L390gat ); 
   BU1 U82 ( L297gat, L391gat ); 
   OR2 U83 ( L270gat, L343gat, L392gat ); 
   IN1 U84 ( L345gat, L393gat ); 
   IN1 U85 ( L346gat, L399gat ); 
   AND2 U86 ( L348gat, L73gat, L400gat ); 
   IN1 U87 ( L349gat, L401gat ); 
   IN1 U88 ( L350gat, L402gat ); 
   IN1 U89 ( L355gat, L403gat ); 
   IN1 U90 ( L357gat, L404gat ); 
   IN1 U91 ( L360gat, L405gat ); 
   AND2 U92 ( L357gat, L360gat, L406gat ); 
   IN1 U93 ( L363gat, L407gat ); 
   IN1 U94 ( L366gat, L408gat ); 
   AND2 U95 ( L363gat, L366gat, L409gat ); 
   NA2 U96 ( L347gat, L352gat, L410gat ); 
   IN1 U97 ( L376gat, L411gat ); 
   IN1 U98 ( L379gat, L412gat ); 
   AND2 U99 ( L376gat, L379gat, L413gat ); 
   IN1 U100 ( L382gat, L414gat ); 
   IN1 U101 ( L385gat, L415gat ); 
   AND2 U102 ( L382gat, L385gat, L416gat ); 
   AND2 U103 ( L210gat, L369gat, L417gat ); 
   BU1 U104 ( L342gat, L418gat ); 
   BU1 U105 ( L344gat, L419gat ); 
   BU1 U106 ( L351gat, L420gat ); 
   BU1 U107 ( L353gat, L421gat ); 
   BU1 U108 ( L354gat, L422gat ); 
   BU1 U109 ( L356gat, L423gat ); 
   IN1 U110 ( L400gat, L424gat ); 
   AND2 U111 ( L404gat, L405gat, L425gat ); 
   AND2 U112 ( L407gat, L408gat, L426gat ); 
   AND3 U113 ( L319gat, L393gat, L55gat, L427gat ); 
   AND3 U114 ( L393gat, L17gat, L287gat, L432gat ); 
   NA3 U115 ( L393gat, L287gat, L55gat, L437gat ); 
   NA4 U116 ( L375gat, L59gat, L156gat, L393gat, L442gat ); 
   NA3 U117 ( L393gat, L319gat, L17gat, L443gat ); 
   AND2 U118 ( L411gat, L412gat, L444gat ); 
   AND2 U119 ( L414gat, L415gat, L445gat ); 
   BU1 U120 ( L392gat, L446gat ); 
   BU1 U121 ( L399gat, L447gat ); 
   BU1 U122 ( L401gat, L448gat ); 
   BU1 U123 ( L402gat, L449gat ); 
   BU1 U124 ( L403gat, L450gat ); 
   IN1 U125 ( L424gat, L451gat ); 
   NO2 U126 ( L406gat, L425gat, L460gat ); 
   NO2 U127 ( L409gat, L426gat, L463gat ); 
   NA2 U128 ( L442gat, L410gat, L466gat ); 
   AND2 U129 ( L143gat, L427gat, L475gat ); 
   AND2 U130 ( L310gat, L432gat, L476gat ); 
   AND2 U131 ( L146gat, L427gat, L477gat ); 
   AND2 U132 ( L310gat, L432gat, L478gat ); 
   AND2 U133 ( L149gat, L427gat, L479gat ); 
   AND2 U134 ( L310gat, L432gat, L480gat ); 
   AND2 U135 ( L153gat, L427gat, L481gat ); 
   AND2 U136 ( L310gat, L432gat, L482gat ); 
   NA2 U137 ( L443gat, L1gat, L483gat ); 
   OR2 U138 ( L369gat, L437gat, L488gat ); 
   OR2 U139 ( L369gat, L437gat, L489gat ); 
   OR2 U140 ( L369gat, L437gat, L490gat ); 
   OR2 U141 ( L369gat, L437gat, L491gat ); 
   NO2 U142 ( L413gat, L444gat, L492gat ); 
   NO2 U143 ( L416gat, L445gat, L495gat ); 
   NA2 U144 ( L130gat, L460gat, L498gat ); 
   OR2 U145 ( L130gat, L460gat, L499gat ); 
   NA2 U146 ( L463gat, L135gat, L500gat ); 
   OR2 U147 ( L463gat, L135gat, L501gat ); 
   AND2 U148 ( L91gat, L466gat, L502gat ); 
   NO2 U149 ( L475gat, L476gat, L503gat ); 
   AND2 U150 ( L96gat, L466gat, L504gat ); 
   NO2 U151 ( L477gat, L478gat, L505gat ); 
   AND2 U152 ( L101gat, L466gat, L506gat ); 
   NO2 U153 ( L479gat, L480gat, L507gat ); 
   AND2 U154 ( L106gat, L466gat, L508gat ); 
   NO2 U155 ( L481gat, L482gat, L509gat ); 
   AND2 U156 ( L143gat, L483gat, L510gat ); 
   AND2 U157 ( L111gat, L466gat, L511gat ); 
   AND2 U158 ( L146gat, L483gat, L512gat ); 
   AND2 U159 ( L116gat, L466gat, L513gat ); 
   AND2 U160 ( L149gat, L483gat, L514gat ); 
   AND2 U161 ( L121gat, L466gat, L515gat ); 
   AND2 U162 ( L153gat, L483gat, L516gat ); 
   AND2 U163 ( L126gat, L466gat, L517gat ); 
   NA2 U164 ( L130gat, L492gat, L518gat ); 
   OR2 U165 ( L130gat, L492gat, L519gat ); 
   NA2 U166 ( L495gat, L207gat, L520gat ); 
   OR2 U167 ( L495gat, L207gat, L521gat ); 
   AND2 U168 ( L451gat, L159gat, L522gat ); 
   AND2 U169 ( L451gat, L165gat, L523gat ); 
   AND2 U170 ( L451gat, L171gat, L524gat ); 
   AND2 U171 ( L451gat, L177gat, L525gat ); 
   AND2 U172 ( L451gat, L183gat, L526gat ); 
   NA2 U173 ( L451gat, L189gat, L527gat ); 
   NA2 U174 ( L451gat, L195gat, L528gat ); 
   NA2 U175 ( L451gat, L201gat, L529gat ); 
   NA2 U176 ( L498gat, L499gat, L530gat ); 
   NA2 U177 ( L500gat, L501gat, L533gat ); 
   NO2 U178 ( L309gat, L502gat, L536gat ); 
   NO2 U179 ( L316gat, L504gat, L537gat ); 
   NO2 U180 ( L317gat, L506gat, L538gat ); 
   NO2 U181 ( L318gat, L508gat, L539gat ); 
   NO2 U182 ( L510gat, L511gat, L540gat ); 
   NO2 U183 ( L512gat, L513gat, L541gat ); 
   NO2 U184 ( L514gat, L515gat, L542gat ); 
   NO2 U185 ( L516gat, L517gat, L543gat ); 
   NA2 U186 ( L518gat, L519gat, L544gat ); 
   NA2 U187 ( L520gat, L521gat, L547gat ); 
   IN1 U188 ( L530gat, L550gat ); 
   IN1 U189 ( L533gat, L551gat ); 
   AND2 U190 ( L530gat, L533gat, L552gat ); 
   NA2 U191 ( L536gat, L503gat, L553gat ); 
   NA2 U192 ( L537gat, L505gat, L557gat ); 
   NA2 U193 ( L538gat, L507gat, L561gat ); 
   NA2 U194 ( L539gat, L509gat, L565gat ); 
   NA2 U195 ( L488gat, L540gat, L569gat ); 
   NA2 U196 ( L489gat, L541gat, L573gat ); 
   NA2 U197 ( L490gat, L542gat, L577gat ); 
   NA2 U198 ( L491gat, L543gat, L581gat ); 
   IN1 U199 ( L544gat, L585gat ); 
   IN1 U200 ( L547gat, L586gat ); 
   AND2 U201 ( L544gat, L547gat, L587gat ); 
   AND2 U202 ( L550gat, L551gat, L588gat ); 
   AND2 U203 ( L585gat, L586gat, L589gat ); 
   NA2 U204 ( L553gat, L159gat, L590gat ); 
   OR2 U205 ( L553gat, L159gat, L593gat ); 
   AND2 U206 ( L246gat, L553gat, L596gat ); 
   NA2 U207 ( L557gat, L165gat, L597gat ); 
   OR2 U208 ( L557gat, L165gat, L600gat ); 
   AND2 U209 ( L246gat, L557gat, L605gat ); 
   NA2 U210 ( L561gat, L171gat, L606gat ); 
   OR2 U211 ( L561gat, L171gat, L609gat ); 
   AND2 U212 ( L246gat, L561gat, L615gat ); 
   NA2 U213 ( L565gat, L177gat, L616gat ); 
   OR2 U214 ( L565gat, L177gat, L619gat ); 
   AND2 U215 ( L246gat, L565gat, L624gat ); 
   NA2 U216 ( L569gat, L183gat, L625gat ); 
   OR2 U217 ( L569gat, L183gat, L628gat ); 
   AND2 U218 ( L246gat, L569gat, L631gat ); 
   NA2 U219 ( L573gat, L189gat, L632gat ); 
   OR2 U220 ( L573gat, L189gat, L635gat ); 
   AND2 U221 ( L246gat, L573gat, L640gat ); 
   NA2 U222 ( L577gat, L195gat, L641gat ); 
   OR2 U223 ( L577gat, L195gat, L644gat ); 
   AND2 U224 ( L246gat, L577gat, L650gat ); 
   NA2 U225 ( L581gat, L201gat, L651gat ); 
   OR2 U226 ( L581gat, L201gat, L654gat ); 
   AND2 U227 ( L246gat, L581gat, L659gat ); 
   NO2 U228 ( L552gat, L588gat, L660gat ); 
   NO2 U229 ( L587gat, L589gat, L661gat ); 
   IN1 U230 ( L590gat, L662gat ); 
   AND2 U231 ( L593gat, L590gat, L665gat ); 
   NO2 U232 ( L596gat, L522gat, L669gat ); 
   IN1 U233 ( L597gat, L670gat ); 
   AND2 U234 ( L600gat, L597gat, L673gat ); 
   NO2 U235 ( L605gat, L523gat, L677gat ); 
   IN1 U236 ( L606gat, L678gat ); 
   AND2 U237 ( L609gat, L606gat, L682gat ); 
   NO2 U238 ( L615gat, L524gat, L686gat ); 
   IN1 U239 ( L616gat, L687gat ); 
   AND2 U240 ( L619gat, L616gat, L692gat ); 
   NO2 U241 ( L624gat, L525gat, L696gat ); 
   IN1 U242 ( L625gat, L697gat ); 
   AND2 U243 ( L628gat, L625gat, L700gat ); 
   NO2 U244 ( L631gat, L526gat, L704gat ); 
   IN1 U245 ( L632gat, L705gat ); 
   AND2 U246 ( L635gat, L632gat, L708gat ); 
   NO2 U247 ( L337gat, L640gat, L712gat ); 
   IN1 U248 ( L641gat, L713gat ); 
   AND2 U249 ( L644gat, L641gat, L717gat ); 
   NO2 U250 ( L339gat, L650gat, L721gat ); 
   IN1 U251 ( L651gat, L722gat ); 
   AND2 U252 ( L654gat, L651gat, L727gat ); 
   NO2 U253 ( L341gat, L659gat, L731gat ); 
   NA2 U254 ( L654gat, L261gat, L732gat ); 
   NA3 U255 ( L644gat, L654gat, L261gat, L733gat ); 
   NA4 U256 ( L635gat, L644gat, L654gat, L261gat, L734gat ); 
   IN1 U257 ( L662gat, L735gat ); 
   AND2 U258 ( L228gat, L665gat, L736gat ); 
   AND2 U259 ( L237gat, L662gat, L737gat ); 
   IN1 U260 ( L670gat, L738gat ); 
   AND2 U261 ( L228gat, L673gat, L739gat ); 
   AND2 U262 ( L237gat, L670gat, L740gat ); 
   IN1 U263 ( L678gat, L741gat ); 
   AND2 U264 ( L228gat, L682gat, L742gat ); 
   AND2 U265 ( L237gat, L678gat, L743gat ); 
   IN1 U266 ( L687gat, L744gat ); 
   AND2 U267 ( L228gat, L692gat, L745gat ); 
   AND2 U268 ( L237gat, L687gat, L746gat ); 
   IN1 U269 ( L697gat, L747gat ); 
   AND2 U270 ( L228gat, L700gat, L748gat ); 
   AND2 U271 ( L237gat, L697gat, L749gat ); 
   IN1 U272 ( L705gat, L750gat ); 
   AND2 U273 ( L228gat, L708gat, L751gat ); 
   AND2 U274 ( L237gat, L705gat, L752gat ); 
   IN1 U275 ( L713gat, L753gat ); 
   AND2 U276 ( L228gat, L717gat, L754gat ); 
   AND2 U277 ( L237gat, L713gat, L755gat ); 
   IN1 U278 ( L722gat, L756gat ); 
   NO2 U279 ( L727gat, L261gat, L757gat ); 
   AND2 U280 ( L727gat, L261gat, L758gat ); 
   AND2 U281 ( L228gat, L727gat, L759gat ); 
   AND2 U282 ( L237gat, L722gat, L760gat ); 
   NA2 U283 ( L644gat, L722gat, L761gat ); 
   NA2 U284 ( L635gat, L713gat, L762gat ); 
   NA3 U285 ( L635gat, L644gat, L722gat, L763gat ); 
   NA2 U286 ( L609gat, L687gat, L764gat ); 
   NA2 U287 ( L600gat, L678gat, L765gat ); 
   NA3 U288 ( L600gat, L609gat, L687gat, L766gat ); 
   BU1 U289 ( L660gat, L767gat ); 
   BU1 U290 ( L661gat, L768gat ); 
   NO2 U291 ( L736gat, L737gat, L769gat ); 
   NO2 U292 ( L739gat, L740gat, L770gat ); 
   NO2 U293 ( L742gat, L743gat, L771gat ); 
   NO2 U294 ( L745gat, L746gat, L772gat ); 
   NA4 U295 ( L750gat, L762gat, L763gat, L734gat, L773gat ); 
   NO2 U296 ( L748gat, L749gat, L777gat ); 
   NA3 U297 ( L753gat, L761gat, L733gat, L778gat ); 
   NO2 U298 ( L751gat, L752gat, L781gat ); 
   NA2 U299 ( L756gat, L732gat, L782gat ); 
   NO2 U300 ( L754gat, L755gat, L785gat ); 
   NO2 U301 ( L757gat, L758gat, L786gat ); 
   NO2 U302 ( L759gat, L760gat, L787gat ); 
   NO2 U303 ( L700gat, L773gat, L788gat ); 
   AND2 U304 ( L700gat, L773gat, L789gat ); 
   NO2 U305 ( L708gat, L778gat, L790gat ); 
   AND2 U306 ( L708gat, L778gat, L791gat ); 
   NO2 U307 ( L717gat, L782gat, L792gat ); 
   AND2 U308 ( L717gat, L782gat, L793gat ); 
   AND2 U309 ( L219gat, L786gat, L794gat ); 
   NA2 U310 ( L628gat, L773gat, L795gat ); 
   NA2 U311 ( L795gat, L747gat, L796gat ); 
   NO2 U312 ( L788gat, L789gat, L802gat ); 
   NO2 U313 ( L790gat, L791gat, L803gat ); 
   NO2 U314 ( L792gat, L793gat, L804gat ); 
   NO2 U315 ( L340gat, L794gat, L805gat ); 
   NO2 U316 ( L692gat, L796gat, L806gat ); 
   AND2 U317 ( L692gat, L796gat, L807gat ); 
   AND2 U318 ( L219gat, L802gat, L808gat ); 
   AND2 U319 ( L219gat, L803gat, L809gat ); 
   AND2 U320 ( L219gat, L804gat, L810gat ); 
   NA4 U321 ( L805gat, L787gat, L731gat, L529gat, L811gat ); 
   NA2 U322 ( L619gat, L796gat, L812gat ); 
   NA3 U323 ( L609gat, L619gat, L796gat, L813gat ); 
   NA4 U324 ( L600gat, L609gat, L619gat, L796gat, L814gat ); 
   NA4 U325 ( L738gat, L765gat, L766gat, L814gat, L815gat ); 
   NA3 U326 ( L741gat, L764gat, L813gat, L819gat ); 
   NA2 U327 ( L744gat, L812gat, L822gat ); 
   NO2 U328 ( L806gat, L807gat, L825gat ); 
   NO2 U329 ( L335gat, L808gat, L826gat ); 
   NO2 U330 ( L336gat, L809gat, L827gat ); 
   NO2 U331 ( L338gat, L810gat, L828gat ); 
   IN1 U332 ( L811gat, L829gat ); 
   NO2 U333 ( L665gat, L815gat, L830gat ); 
   AND2 U334 ( L665gat, L815gat, L831gat ); 
   NO2 U335 ( L673gat, L819gat, L832gat ); 
   AND2 U336 ( L673gat, L819gat, L833gat ); 
   NO2 U337 ( L682gat, L822gat, L834gat ); 
   AND2 U338 ( L682gat, L822gat, L835gat ); 
   AND2 U339 ( L219gat, L825gat, L836gat ); 
   NA3 U340 ( L826gat, L777gat, L704gat, L837gat ); 
   NA4 U341 ( L827gat, L781gat, L712gat, L527gat, L838gat ); 
   NA4 U342 ( L828gat, L785gat, L721gat, L528gat, L839gat ); 
   IN1 U343 ( L829gat, L840gat ); 
   NA2 U344 ( L815gat, L593gat, L841gat ); 
   NO2 U345 ( L830gat, L831gat, L842gat ); 
   NO2 U346 ( L832gat, L833gat, L843gat ); 
   NO2 U347 ( L834gat, L835gat, L844gat ); 
   NO2 U348 ( L334gat, L836gat, L845gat ); 
   IN1 U349 ( L837gat, L846gat ); 
   IN1 U350 ( L838gat, L847gat ); 
   IN1 U351 ( L839gat, L848gat ); 
   AND2 U352 ( L735gat, L841gat, L849gat ); 
   BU1 U353 ( L840gat, L850gat ); 
   AND2 U354 ( L219gat, L842gat, L851gat ); 
   AND2 U355 ( L219gat, L843gat, L852gat ); 
   AND2 U356 ( L219gat, L844gat, L853gat ); 
   NA3 U357 ( L845gat, L772gat, L696gat, L854gat ); 
   IN1 U358 ( L846gat, L855gat ); 
   IN1 U359 ( L847gat, L856gat ); 
   IN1 U360 ( L848gat, L857gat ); 
   IN1 U361 ( L849gat, L858gat ); 
   NO2 U362 ( L417gat, L851gat, L859gat ); 
   NO2 U363 ( L332gat, L852gat, L860gat ); 
   NO2 U364 ( L333gat, L853gat, L861gat ); 
   IN1 U365 ( L854gat, L862gat ); 
   BU1 U366 ( L855gat, L863gat ); 
   BU1 U367 ( L856gat, L864gat ); 
   BU1 U368 ( L857gat, L865gat ); 
   BU1 U369 ( L858gat, L866gat ); 
   NA3 U370 ( L859gat, L769gat, L669gat, L867gat ); 
   NA3 U371 ( L860gat, L770gat, L677gat, L868gat ); 
   NA3 U372 ( L861gat, L771gat, L686gat, L869gat ); 
   IN1 U373 ( L862gat, L870gat ); 
   IN1 U374 ( L867gat, L871gat ); 
   IN1 U375 ( L868gat, L872gat ); 
   IN1 U376 ( L869gat, L873gat ); 
   BU1 U377 ( L870gat, L874gat ); 
   IN1 U378 ( L871gat, L875gat ); 
   IN1 U379 ( L872gat, L876gat ); 
   IN1 U380 ( L873gat, L877gat ); 
   BU1 U381 ( L875gat, L878gat ); 
   BU1 U382 ( L876gat, L879gat ); 
   BU1 U383 ( L877gat, L880gat ); 
endmodule

