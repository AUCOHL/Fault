
module c880g ( L1gat, L8gat, L13gat, L17gat, L26gat, L29gat, L36gat, L42gat, 
    L51gat, L55gat, L59gat, L68gat, L72gat, L73gat, L74gat, L75gat, L80gat, 
    L85gat, L86gat, L87gat, L88gat, L89gat, L90gat, L91gat, L96gat, L101gat, 
    L106gat, L111gat, L116gat, L121gat, L126gat, L130gat, L135gat, L138gat, 
    L143gat, L146gat, L149gat, L152gat, L153gat, L156gat, L159gat, L165gat, 
    L171gat, L177gat, L183gat, L189gat, L195gat, L201gat, L207gat, L210gat, 
    L219gat, L228gat, L237gat, L246gat, L255gat, L259gat, L260gat, L261gat, 
    L267gat, L268gat, L388gat, L389gat, L390gat, L391gat, L418gat, L419gat, 
    L420gat, L421gat, L422gat, L423gat, L446gat, L447gat, L448gat, L449gat, 
    L450gat, L767gat, L768gat, L850gat, L863gat, L864gat, L865gat, L866gat, 
    L874gat, L878gat, L879gat, L880gat );
input  L1gat, L8gat, L13gat, L17gat, L26gat, L29gat, L36gat, L42gat, L51gat, 
    L55gat, L59gat, L68gat, L72gat, L73gat, L74gat, L75gat, L80gat, L85gat, 
    L86gat, L87gat, L88gat, L89gat, L90gat, L91gat, L96gat, L101gat, L106gat, 
    L111gat, L116gat, L121gat, L126gat, L130gat, L135gat, L138gat, L143gat, 
    L146gat, L149gat, L152gat, L153gat, L156gat, L159gat, L165gat, L171gat, 
    L177gat, L183gat, L189gat, L195gat, L201gat, L207gat, L210gat, L219gat, 
    L228gat, L237gat, L246gat, L255gat, L259gat, L260gat, L261gat, L267gat, 
    L268gat;
output L388gat, L389gat, L390gat, L391gat, L418gat, L419gat, L420gat, L421gat, 
    L422gat, L423gat, L446gat, L447gat, L448gat, L449gat, L450gat, L767gat, 
    L768gat, L850gat, L863gat, L864gat, L865gat, L866gat, L874gat, L878gat, 
    L879gat, L880gat;
    tri L1gat_wire, L269gat, L29gat_wire, L87gat_wire, L165gat_wire, 
        L446gat_wire, L759gat, L804gat, L529gat, L587gat, L391gat_wire, 
        L876gat, L503gat, L644gat, L773gat, L785gat, L880gat_wire, L303gat, 
        L306gat, L625gat, L712gat, L382gat, L427gat, L489gat, L510gat, L738gat, 
        L796gat, L865gat_wire, L678gat, L760gat, L450gat_wire, L717gat, 
        L812gat, L74gat_wire, L91gat_wire, L329gat, L408gat, L101gat_wire, 
        L765gat, L860gat, L138gat_wire, L310gat, L159gat_wire, L422gat_wire, 
        L515gat, L246gat_wire, L793gat, L348gat, L838gat, L704gat, L443gat, 
        L619gat, L859gat, L152gat_wire, L255gat_wire, L506gat, L641gat, 
        L736gat, L873gat, L833gat, L322gat, L267gat_wire, L659gat, L819gat, 
        L350gat, L403gat, L744gat, L8gat_wire, L26gat_wire, L55gat_wire, 
        L291gat, L673gat, L841gat, L308gat, L331gat, L878gat_wire, L343gat, 
        L89gat_wire, L369gat, L448gat_wire, L660gat, L757gat, L852gat, L410gat, 
        L696gat, L527gat, L589gat, L287gat, L334gat, L491gat, L508gat, L825gat, 
        L550gat, L346gat, L415gat, L778gat, L522gat, L857gat, L290gat, L294gat, 
        L327gat, L389gat_wire, L665gat, L752gat, L543gat, L210gat_wire, 
        L482gat, L836gat, L569gat, L733gat, L844gat, L351gat, L355gat, L406gat, 
        L741gat, L402gat, L121gat_wire, L840gat, L309gat, L745gat, L323gat, 
        L153gat_wire, L832gat, L547gat, L600gat, L737gat, L342gat, L411gat, 
        L449gat_wire, L526gat, L661gat, L853gat, L756gat, L697gat, L588gat, 
        L879gat_wire, L270gat, L51gat_wire, L88gat_wire, L330gat, L463gat, 
        L207gat_wire, L495gat, L347gat, L36gat_wire, L42gat_wire, L286gat, 
        L414gat, L523gat, L692gat, L753gat, L295gat, L335gat, L490gat, L509gat, 
        L228gat_wire, L856gat, L721gat, L616gat, L466gat, L551gat, L677gat, 
        L740gat, L354gat, L845gat, L407gat, L530gat, L276gat, L280gat, 
        L68gat_wire, L326gat, L388gat_wire, L475gat, L542gat, L732gat, 
        L75gat_wire, L86gat_wire, L156gat_wire, L483gat, L605gat, L837gat, 
        L302gat, L116gat_wire, L390gat_wire, L772gat, L877gat, L307gat, 
        L268gat_wire, L366gat, L375gat, L447gat_wire, L502gat, L758gat, 
        L488gat, L528gat, L586gat, L700gat, L805gat, L739gat, L426gat, L511gat, 
        L761gat, L864gat_wire, L177gat_wire, L624gat, L713gat, L328gat, 
        L90gat_wire, L423gat_wire, L764gat, L861gat, L451gat, L514gat, L792gat, 
        L839gat, L409gat, L590gat, L813gat, L333gat, L349gat, L363gat, L507gat, 
        L781gat, L640gat, L777gat, L872gat, L442gat, L632gat, L705gat, L460gat, 
        L557gat, L858gat, L143gat_wire, L789gat, L822gat, L727gat, 
        L850gat_wire, L319gat, L662gat, L755gat, L412gat, L808gat, L525gat, 
        L341gat, L734gat, L831gat, L869gat, L352gat, L401gat, L544gat, L687gat, 
        L536gat, L13gat_wire, L17gat_wire, L273gat, L293gat, L843gat, L296gat, 
        L325gat, L746gat, L476gat, L541gat, L480gat, L519gat, L769gat, L606gat, 
        L731gat, L743gat, L834gat, L846gat, L189gat_wire, L201gat_wire, 
        L336gat, L259gat_wire, L260gat_wire, L357gat, L404gat, L682gat, 
        L146gat_wire, L533gat, L615gat, L722gat, L827gat, L552gat, L59gat_wire, 
        L285gat, L344gat, L417gat, L520gat, L708gat, L750gat, L855gat, 
        L96gat_wire, L304gat, L538gat, L596gat, L815gat, L748gat, L376gat, 
        L425gat, L512gat, L794gat, L219gat_wire, L106gat_wire, L762gat, 
        L867gat, L317gat, L444gat, L573gat, L585gat, L80gat_wire, L85gat_wire, 
        L393gat, L771gat, L806gat, L874gat_wire, L360gat, L73gat_wire, 
        L419gat_wire, L498gat, L501gat, L631gat, L787gat, L803gat, L504gat, 
        L669gat, L782gat, L829gat, L298gat, L301gat, L338gat, L565gat, L871gat, 
        L848gat, L171gat_wire, L810gat, L385gat, L593gat, L420gat_wire, 
        L478gat, L650gat, L862gat, L767gat_wire, L517gat, L791gat, L424gat, 
        L513gat, L539gat, L597gat, L654gat, L763gat, L795gat, L866gat_wire, 
        L814gat, L279gat, L72gat_wire, L305gat, L183gat_wire, L561gat, L749gat, 
        L392gat, L875gat, L770gat, L316gat, L437gat, L499gat, L445gat, L500gat, 
        L786gat, L284gat, L292gat, L111gat_wire, L339gat, L432gat, L635gat, 
        L807gat, L149gat_wire, L505gat, L828gat, L870gat, L318gat, 
        L195gat_wire, L418gat_wire, L581gat, L802gat, L421gat_wire, L479gat, 
        L577gat, L651gat, L766gat, L863gat_wire, L609gat, L130gat_wire, 
        L516gat, L237gat_wire, L790gat, L754gat, L811gat, L849gat, L851gat, 
        L332gat, L340gat, L809gat, L413gat, L524gat, L353gat, L788gat, L400gat, 
        L537gat, L686gat, L628gat, L670gat, L747gat, L297gat, L379gat, L735gat, 
        L842gat, L830gat, L868gat, L126gat_wire, L847gat, L324gat, L356gat, 
        L405gat, L742gat, L477gat, L261gat_wire, L540gat, L345gat, L416gat, 
        L481gat, L518gat, L768gat_wire, L835gat, L521gat, L337gat, L399gat, 
        L492gat, L135gat_wire, L854gat, L751gat, L826gat, L553gat;
    assign L1gat_wire = L1gat;
    assign L8gat_wire = L8gat;
    assign L13gat_wire = L13gat;
    assign L17gat_wire = L17gat;
    assign L26gat_wire = L26gat;
    assign L29gat_wire = L29gat;
    assign L36gat_wire = L36gat;
    assign L42gat_wire = L42gat;
    assign L51gat_wire = L51gat;
    assign L55gat_wire = L55gat;
    assign L59gat_wire = L59gat;
    assign L68gat_wire = L68gat;
    assign L72gat_wire = L72gat;
    assign L73gat_wire = L73gat;
    assign L74gat_wire = L74gat;
    assign L75gat_wire = L75gat;
    assign L80gat_wire = L80gat;
    assign L85gat_wire = L85gat;
    assign L86gat_wire = L86gat;
    assign L87gat_wire = L87gat;
    assign L88gat_wire = L88gat;
    assign L89gat_wire = L89gat;
    assign L90gat_wire = L90gat;
    assign L91gat_wire = L91gat;
    assign L96gat_wire = L96gat;
    assign L101gat_wire = L101gat;
    assign L106gat_wire = L106gat;
    assign L111gat_wire = L111gat;
    assign L116gat_wire = L116gat;
    assign L121gat_wire = L121gat;
    assign L126gat_wire = L126gat;
    assign L130gat_wire = L130gat;
    assign L135gat_wire = L135gat;
    assign L138gat_wire = L138gat;
    assign L143gat_wire = L143gat;
    assign L146gat_wire = L146gat;
    assign L149gat_wire = L149gat;
    assign L152gat_wire = L152gat;
    assign L153gat_wire = L153gat;
    assign L156gat_wire = L156gat;
    assign L159gat_wire = L159gat;
    assign L165gat_wire = L165gat;
    assign L171gat_wire = L171gat;
    assign L177gat_wire = L177gat;
    assign L183gat_wire = L183gat;
    assign L189gat_wire = L189gat;
    assign L195gat_wire = L195gat;
    assign L201gat_wire = L201gat;
    assign L207gat_wire = L207gat;
    assign L210gat_wire = L210gat;
    assign L219gat_wire = L219gat;
    assign L228gat_wire = L228gat;
    assign L237gat_wire = L237gat;
    assign L246gat_wire = L246gat;
    assign L255gat_wire = L255gat;
    assign L259gat_wire = L259gat;
    assign L260gat_wire = L260gat;
    assign L261gat_wire = L261gat;
    assign L267gat_wire = L267gat;
    assign L268gat_wire = L268gat;
    assign L388gat = L388gat_wire;
    assign L389gat = L389gat_wire;
    assign L390gat = L390gat_wire;
    assign L391gat = L391gat_wire;
    assign L418gat = L418gat_wire;
    assign L419gat = L419gat_wire;
    assign L420gat = L420gat_wire;
    assign L421gat = L421gat_wire;
    assign L422gat = L422gat_wire;
    assign L423gat = L423gat_wire;
    assign L446gat = L446gat_wire;
    assign L447gat = L447gat_wire;
    assign L448gat = L448gat_wire;
    assign L449gat = L449gat_wire;
    assign L450gat = L450gat_wire;
    assign L767gat = L767gat_wire;
    assign L768gat = L768gat_wire;
    assign L850gat = L850gat_wire;
    assign L863gat = L863gat_wire;
    assign L864gat = L864gat_wire;
    assign L865gat = L865gat_wire;
    assign L866gat = L866gat_wire;
    assign L874gat = L874gat_wire;
    assign L878gat = L878gat_wire;
    assign L879gat = L879gat_wire;
    assign L880gat = L880gat_wire;
    nand4 U1 ( L1gat_wire, L8gat_wire, L13gat_wire, L17gat_wire, L269gat );
    nand4 U6 ( L1gat_wire, L8gat_wire, L13gat_wire, L55gat_wire, L280gat );
    and3 U14 ( L59gat_wire, L75gat_wire, L80gat_wire, L293gat );
    or2 U21 ( L91gat_wire, L96gat_wire, L302gat );
    inv U54 ( L269gat, L342gat );
    inv U73 ( L310gat, L369gat );
    and3 U113 ( L319gat, L393gat, L55gat_wire, L427gat );
    or2 U223 ( L577gat, L195gat_wire, L644gat );
    and2 U134 ( L310gat, L432gat, L480gat );
    nand2 U96 ( L347gat, L352gat, L410gat );
    nand2 U198 ( L491gat, L543gat, L581gat );
    nand2 U204 ( L553gat, L159gat_wire, L590gat );
    and2 U338 ( L682gat, L822gat, L835gat );
    and2 U356 ( L219gat_wire, L844gat, L853gat );
    nand3 U371 ( L860gat, L770gat, L677gat, L868gat );
    nand2 U166 ( L495gat, L207gat_wire, L520gat );
    nand4 U256 ( L635gat, L644gat, L654gat, L261gat_wire, L734gat );
    and2 U271 ( L237gat_wire, L697gat, L749gat );
    and2 U68 ( L90gat_wire, L298gat, L356gat );
    buffer U108 ( L354gat, L422gat_wire );
    or2 U141 ( L369gat, L437gat, L491gat );
    nor2 U183 ( L512gat, L513gat, L541gat );
    nor2 U294 ( L745gat, L746gat, L772gat );
    and2 U304 ( L700gat, L773gat, L789gat );
    nand3 U323 ( L609gat, L619gat, L796gat, L813gat );
    nor2 U238 ( L615gat, L524gat, L686gat );
    nand2 U174 ( L451gat, L195gat_wire, L528gat );
    nand2 U191 ( L536gat, L503gat, L553gat );
    nand2 U286 ( L609gat, L687gat, L764gat );
    nor2 U316 ( L692gat, L796gat, L806gat );
    nor2 U331 ( L338gat, L810gat, L828gat );
    inv U378 ( L871gat, L875gat );
    nor2 U244 ( L631gat, L526gat, L704gat );
    and2 U28 ( L8gat_wire, L138gat_wire, L309gat );
    nand2 U33 ( L59gat_wire, L156gat_wire, L319gat );
    inv U263 ( L678gat, L741gat );
    and2 U148 ( L91gat_wire, L466gat, L502gat );
    nor2 U153 ( L479gat, L480gat, L507gat );
    inv U278 ( L722gat, L756gat );
    or2 U41 ( L183gat_wire, L189gat_wire, L329gat );
    and2 U46 ( L210gat_wire, L101gat_wire, L334gat );
    or2 U61 ( L280gat, L285gat, L349gat );
    inv U84 ( L345gat, L393gat );
    nand2 U344 ( L815gat, L593gat, L841gat );
    nor2 U363 ( L332gat, L852gat, L860gat );
    inv U101 ( L385gat, L415gat );
    and2 U231 ( L593gat, L590gat, L665gat );
    nor2 U126 ( L406gat, L425gat, L460gat );
    or2 U211 ( L561gat, L171gat_wire, L609gat );
    nand2 U216 ( L569gat, L183gat_wire, L625gat );
    buffer U381 ( L875gat, L878gat_wire );
    inv U66 ( L296gat, L354gat );
    buffer U106 ( L351gat, L420gat_wire );
    buffer U121 ( L399gat, L447gat_wire );
    inv U236 ( L606gat, L678gat );
    and2 U168 ( L451gat, L159gat_wire, L522gat );
    nand4 U2 ( L1gat_wire, L26gat_wire, L13gat_wire, L17gat_wire, L270gat );
    nand4 U5 ( L1gat_wire, L8gat_wire, L51gat_wire, L17gat_wire, L279gat );
    nand4 U7 ( L59gat_wire, L42gat_wire, L68gat_wire, L72gat_wire, L284gat );
    nand2 U8 ( L29gat_wire, L68gat_wire, L285gat );
    and3 U13 ( L29gat_wire, L36gat_wire, L42gat_wire, L292gat );
    nor2 U34 ( L17gat_wire, L42gat_wire, L322gat );
    or2 U83 ( L270gat, L343gat, L392gat );
    and2 U258 ( L228gat_wire, L665gat, L736gat );
    inv U98 ( L379gat, L412gat );
    inv U343 ( L829gat, L840gat );
    inv U358 ( L846gat, L855gat );
    nor2 U364 ( L333gat, L853gat, L861gat );
    and2 U154 ( L106gat_wire, L466gat, L508gat );
    and2 U264 ( L228gat_wire, L682gat, L742gat );
    nand2 U26 ( L121gat_wire, L126gat_wire, L307gat );
    and2 U48 ( L210gat_wire, L111gat_wire, L336gat );
    nand2 U128 ( L442gat, L410gat, L466gat );
    nand2 U173 ( L451gat, L189gat_wire, L527gat );
    and2 U243 ( L628gat, L625gat, L700gat );
    nor2 U184 ( L514gat, L515gat, L542gat );
    nand2 U196 ( L489gat, L541gat, L573gat );
    and2 U336 ( L673gat, L819gat, L833gat );
    and2 U281 ( L228gat_wire, L727gat, L759gat );
    nand2 U311 ( L795gat, L747gat, L796gat );
    nand4 U324 ( L600gat, L609gat, L619gat, L796gat, L814gat );
    nor2 U293 ( L742gat, L743gat, L771gat );
    nor2 U303 ( L700gat, L773gat, L788gat );
    nand2 U146 ( L463gat, L135gat_wire, L500gat );
    and2 U218 ( L246gat_wire, L569gat, L631gat );
    inv U251 ( L651gat, L722gat );
    and2 U276 ( L228gat_wire, L717gat, L754gat );
    nand3 U9 ( L59gat_wire, L68gat_wire, L74gat_wire, L286gat );
    and3 U12 ( L29gat_wire, L36gat_wire, L80gat_wire, L291gat );
    and2 U35 ( L17gat_wire, L42gat_wire, L323gat );
    and2 U53 ( L255gat_wire, L267gat_wire, L341gat );
    inv U91 ( L360gat, L405gat );
    and2 U161 ( L121gat_wire, L466gat, L515gat );
    and2 U203 ( L585gat, L586gat, L589gat );
    inv U351 ( L839gat, L848gat );
    inv U376 ( L869gat, L873gat );
    nor2 U74 ( L322gat, L323gat, L375gat );
    and3 U114 ( L393gat, L17gat_wire, L287gat, L432gat );
    and2 U133 ( L149gat_wire, L427gat, L479gat );
    and2 U224 ( L246gat_wire, L577gat, L650gat );
    and2 U99 ( L376gat, L379gat, L413gat );
    nand2 U197 ( L490gat, L542gat, L577gat );
    nand3 U288 ( L600gat, L609gat, L687gat, L766gat );
    and2 U318 ( L219gat_wire, L802gat, L808gat );
    nor2 U337 ( L682gat, L822gat, L834gat );
    and2 U280 ( L727gat, L261gat_wire, L758gat );
    nand2 U310 ( L628gat, L773gat, L795gat );
    nor2 U155 ( L481gat, L482gat, L509gat );
    inv U359 ( L847gat, L856gat );
    and2 U265 ( L237gat_wire, L678gat, L743gat );
    inv U242 ( L625gat, L697gat );
    or2 U27 ( L121gat_wire, L126gat_wire, L308gat );
    nand2 U40 ( L183gat_wire, L189gat_wire, L328gat );
    buffer U82 ( L297gat, L391gat_wire );
    and2 U169 ( L451gat, L165gat_wire, L523gat );
    and2 U172 ( L451gat, L183gat_wire, L526gat );
    and2 U259 ( L237gat_wire, L662gat, L737gat );
    nand4 U342 ( L828gat, L785gat, L721gat, L528gat, L839gat );
    inv U365 ( L854gat, L862gat );
    and2 U52 ( L210gat_wire, L121gat_wire, L340gat );
    nand2 U67 ( L89gat_wire, L298gat, L355gat );
    buffer U107 ( L353gat, L421gat_wire );
    buffer U120 ( L392gat, L446gat_wire );
    nand2 U210 ( L561gat, L171gat_wire, L606gat );
    inv U380 ( L873gat, L877gat );
    and2 U237 ( L609gat, L606gat, L682gat );
    nand2 U75 ( L324gat, L325gat, L376gat );
    nand3 U115 ( L393gat, L287gat, L55gat_wire, L437gat );
    and2 U132 ( L310gat, L432gat, L478gat );
    and2 U202 ( L550gat, L551gat, L588gat );
    inv U90 ( L357gat, L404gat );
    nand2 U225 ( L581gat, L201gat_wire, L651gat );
    buffer U289 ( L660gat, L767gat_wire );
    and2 U319 ( L219gat_wire, L803gat, L809gat );
    inv U350 ( L838gat, L847gat );
    or2 U147 ( L463gat, L135gat_wire, L501gat );
    buffer U377 ( L870gat, L874gat_wire );
    and2 U277 ( L237gat_wire, L713gat, L755gat );
    and2 U160 ( L149gat_wire, L483gat, L514gat );
    nor2 U250 ( L339gat, L650gat, L721gat );
    nand2 U20 ( L91gat_wire, L96gat_wire, L301gat );
    and2 U49 ( L255gat_wire, L259gat_wire, L337gat );
    and2 U129 ( L143gat_wire, L427gat, L475gat );
    nor2 U185 ( L516gat, L517gat, L543gat );
    nand4 U325 ( L738gat, L765gat, L766gat, L814gat, L815gat );
    nor2 U292 ( L739gat, L740gat, L770gat );
    nor2 U302 ( L759gat, L760gat, L787gat );
    nand2 U219 ( L573gat, L189gat_wire, L632gat );
    nand2 U69 ( L301gat, L302gat, L357gat );
    buffer U109 ( L356gat, L423gat_wire );
    nor2 U182 ( L510gat, L511gat, L540gat );
    nand4 U295 ( L750gat, L762gat, L763gat, L734gat, L773gat );
    nor2 U305 ( L708gat, L778gat, L790gat );
    nand2 U322 ( L619gat, L796gat, L812gat );
    or2 U167 ( L495gat, L207gat_wire, L521gat );
    inv U239 ( L616gat, L687gat );
    inv U257 ( L662gat, L735gat );
    inv U29 ( L268gat_wire, L310gat );
    and2 U47 ( L210gat_wire, L106gat_wire, L335gat );
    inv U55 ( L273gat, L343gat );
    nand2 U72 ( L307gat, L308gat, L366gat );
    inv U97 ( L376gat, L411gat );
    or2 U140 ( L369gat, L437gat, L490gat );
    and2 U270 ( L228gat_wire, L700gat, L748gat );
    nand3 U370 ( L859gat, L769gat, L669gat, L867gat );
    nand2 U222 ( L577gat, L195gat_wire, L641gat );
    nand3 U357 ( L845gat, L772gat, L696gat, L854gat );
    and2 U112 ( L407gat, L408gat, L426gat );
    and2 U135 ( L153gat_wire, L427gat, L481gat );
    or2 U205 ( L553gat, L159gat_wire, L593gat );
    nor2 U60 ( L280gat, L284gat, L348gat );
    inv U199 ( L544gat, L585gat );
    and2 U339 ( L219gat_wire, L825gat, L836gat );
    inv U230 ( L590gat, L662gat );
    inv U100 ( L382gat, L414gat );
    nor2 U127 ( L409gat, L426gat, L463gat );
    or2 U217 ( L569gat, L183gat_wire, L628gat );
    nor2 U149 ( L475gat, L476gat, L503gat );
    nor2 U279 ( L727gat, L261gat_wire, L757gat );
    and3 U15 ( L59gat_wire, L75gat_wire, L42gat_wire, L294gat );
    inv U85 ( L346gat, L399gat );
    nor2 U362 ( L417gat, L851gat, L859gat );
    nand2 U175 ( L451gat, L201gat_wire, L529gat );
    nor2 U345 ( L830gat, L831gat, L842gat );
    inv U379 ( L872gat, L876gat );
    and3 U17 ( L59gat_wire, L36gat_wire, L42gat_wire, L296gat );
    nand2 U22 ( L101gat_wire, L106gat_wire, L303gat );
    and2 U32 ( L152gat_wire, L138gat_wire, L318gat );
    inv U245 ( L632gat, L705gat );
    or2 U39 ( L171gat_wire, L177gat_wire, L327gat );
    inv U57 ( L276gat, L345gat );
    nand2 U137 ( L443gat, L1gat_wire, L483gat );
    and2 U152 ( L101gat_wire, L466gat, L506gat );
    and2 U262 ( L237gat_wire, L670gat, L740gat );
    and2 U190 ( L530gat, L533gat, L552gat );
    nand2 U287 ( L600gat, L678gat, L765gat );
    and2 U317 ( L692gat, L796gat, L807gat );
    nor2 U330 ( L336gat, L809gat, L827gat );
    nand2 U70 ( L303gat, L304gat, L360gat );
    nand2 U207 ( L557gat, L165gat_wire, L597gat );
    inv U110 ( L400gat, L424gat );
    or2 U220 ( L573gat, L189gat_wire, L635gat );
    and2 U159 ( L116gat_wire, L466gat, L513gat );
    and2 U95 ( L363gat, L366gat, L409gat );
    inv U269 ( L697gat, L747gat );
    and2 U355 ( L219gat_wire, L843gat, L852gat );
    inv U272 ( L705gat, L750gat );
    buffer U369 ( L858gat, L866gat_wire );
    nand3 U372 ( L861gat, L771gat, L686gat, L869gat );
    and2 U30 ( L51gat_wire, L138gat_wire, L316gat );
    buffer U79 ( L290gat, L388gat_wire );
    and2 U119 ( L414gat, L415gat, L445gat );
    nor2 U142 ( L413gat, L444gat, L492gat );
    or2 U165 ( L130gat_wire, L492gat, L519gat );
    nor2 U180 ( L317gat, L506gat, L538gat );
    nand3 U255 ( L644gat, L654gat, L261gat_wire, L733gat );
    nand2 U192 ( L537gat, L505gat, L557gat );
    nand3 U297 ( L753gat, L761gat, L733gat, L778gat );
    and2 U320 ( L219gat_wire, L804gat, L810gat );
    nor2 U307 ( L717gat, L782gat, L792gat );
    nand3 U285 ( L635gat, L644gat, L722gat, L763gat );
    nor2 U315 ( L340gat, L794gat, L805gat );
    inv U332 ( L811gat, L829gat );
    nor2 U229 ( L587gat, L589gat, L661gat );
    inv U260 ( L670gat, L738gat );
    and2 U150 ( L96gat_wire, L466gat, L504gat );
    nand2 U177 ( L500gat, L501gat, L533gat );
    nor2 U247 ( L337gat, L640gat, L712gat );
    inv U87 ( L349gat, L401gat );
    nor2 U347 ( L834gat, L835gat, L844gat );
    inv U360 ( L848gat, L857gat );
    nand2 U42 ( L195gat_wire, L201gat_wire, L330gat );
    and2 U45 ( L210gat_wire, L96gat_wire, L333gat );
    inv U125 ( L424gat, L451gat );
    or2 U62 ( L280gat, L286gat, L350gat );
    and2 U215 ( L246gat_wire, L565gat, L624gat );
    inv U65 ( L295gat, L353gat );
    and2 U102 ( L382gat, L385gat, L416gat );
    nor2 U232 ( L596gat, L522gat, L669gat );
    buffer U105 ( L344gat, L419gat_wire );
    inv U189 ( L533gat, L551gat );
    nor2 U329 ( L335gat, L808gat, L826gat );
    nor2 U235 ( L605gat, L523gat, L677gat );
    and2 U212 ( L246gat_wire, L561gat, L615gat );
    buffer U382 ( L876gat, L879gat_wire );
    buffer U80 ( L291gat, L389gat_wire );
    buffer U122 ( L401gat, L448gat_wire );
    nand2 U299 ( L756gat, L732gat, L782gat );
    and2 U309 ( L219gat_wire, L786gat, L794gat );
    buffer U367 ( L856gat, L864gat_wire );
    nand3 U340 ( L826gat, L777gat, L704gat, L837gat );
    and3 U3 ( L29gat_wire, L36gat_wire, L42gat_wire, L273gat );
    and3 U10 ( L29gat_wire, L75gat_wire, L80gat_wire, L287gat );
    and3 U11 ( L29gat_wire, L75gat_wire, L42gat_wire, L290gat );
    or2 U19 ( L87gat_wire, L88gat_wire, L298gat );
    or2 U25 ( L111gat_wire, L116gat_wire, L306gat );
    or2 U37 ( L159gat_wire, L165gat_wire, L325gat );
    and2 U157 ( L111gat_wire, L466gat, L511gat );
    and2 U170 ( L451gat, L171gat_wire, L524gat );
    and2 U240 ( L619gat, L616gat, L692gat );
    inv U59 ( L279gat, L347gat );
    or2 U139 ( L369gat, L437gat, L489gat );
    nand2 U195 ( L488gat, L540gat, L569gat );
    and2 U267 ( L228gat_wire, L692gat, L745gat );
    and2 U282 ( L237gat_wire, L722gat, L760gat );
    nor2 U312 ( L788gat, L789gat, L802gat );
    nor2 U335 ( L673gat, L819gat, L832gat );
    inv U89 ( L355gat, L403gat );
    nand2 U187 ( L520gat, L521gat, L547gat );
    and2 U209 ( L246gat_wire, L557gat, L605gat );
    buffer U290 ( L661gat, L768gat_wire );
    nor2 U300 ( L754gat, L755gat, L785gat );
    nand2 U327 ( L744gat, L812gat, L822gat );
    inv U349 ( L837gat, L846gat );
    or2 U145 ( L130gat_wire, L460gat, L499gat );
    and2 U162 ( L153gat_wire, L483gat, L516gat );
    and2 U252 ( L654gat, L651gat, L727gat );
    nor2 U179 ( L316gat, L504gat, L537gat );
    inv U275 ( L713gat, L753gat );
    and2 U249 ( L644gat, L641gat, L717gat );
    and2 U50 ( L210gat_wire, L116gat_wire, L338gat );
    nand2 U77 ( L328gat, L329gat, L382gat );
    and2 U92 ( L357gat, L360gat, L406gat );
    inv U375 ( L868gat, L872gat );
    nand3 U117 ( L393gat, L319gat, L17gat_wire, L443gat );
    and2 U352 ( L735gat, L841gat, L849gat );
    and2 U227 ( L246gat_wire, L581gat, L659gat );
    inv U200 ( L547gat, L586gat );
    inv U58 ( L276gat, L346gat );
    and2 U130 ( L310gat, L432gat, L476gat );
    or2 U138 ( L369gat, L437gat, L488gat );
    nand2 U194 ( L539gat, L509gat, L565gat );
    nand2 U283 ( L644gat, L722gat, L761gat );
    nor2 U313 ( L790gat, L791gat, L803gat );
    and2 U334 ( L665gat, L815gat, L831gat );
    or2 U208 ( L557gat, L165gat_wire, L600gat );
    nor2 U241 ( L624gat, L525gat, L696gat );
    nand2 U36 ( L159gat_wire, L165gat_wire, L324gat );
    and2 U156 ( L143gat_wire, L483gat, L510gat );
    and2 U171 ( L451gat, L177gat_wire, L525gat );
    inv U266 ( L687gat, L744gat );
    buffer U81 ( L292gat, L390gat_wire );
    nand4 U341 ( L827gat, L781gat, L712gat, L527gat, L838gat );
    buffer U366 ( L855gat, L863gat_wire );
    and3 U4 ( L1gat_wire, L26gat_wire, L51gat_wire, L276gat );
    and2 U18 ( L85gat_wire, L86gat_wire, L297gat );
    or2 U43 ( L195gat_wire, L201gat_wire, L331gat );
    inv U64 ( L294gat, L352gat );
    buffer U104 ( L342gat, L418gat_wire );
    and2 U234 ( L600gat, L597gat, L673gat );
    and2 U51 ( L255gat_wire, L260gat_wire, L339gat );
    nand2 U76 ( L326gat, L327gat, L379gat );
    nand4 U116 ( L375gat, L59gat_wire, L156gat_wire, L393gat, L442gat );
    buffer U123 ( L402gat, L449gat_wire );
    nand2 U213 ( L565gat, L177gat_wire, L616gat );
    buffer U383 ( L877gat, L880gat_wire );
    nor2 U298 ( L751gat, L752gat, L781gat );
    and2 U308 ( L717gat, L782gat, L793gat );
    or2 U226 ( L581gat, L201gat_wire, L654gat );
    and2 U131 ( L146gat_wire, L427gat, L477gat );
    and2 U201 ( L544gat, L547gat, L587gat );
    nor2 U178 ( L309gat, L502gat, L536gat );
    or2 U23 ( L101gat_wire, L106gat_wire, L304gat );
    nand2 U24 ( L111gat_wire, L116gat_wire, L305gat );
    inv U88 ( L350gat, L402gat );
    inv U93 ( L363gat, L407gat );
    inv U248 ( L641gat, L713gat );
    buffer U353 ( L840gat, L850gat_wire );
    inv U374 ( L867gat, L871gat );
    nand2 U144 ( L130gat_wire, L460gat, L498gat );
    and2 U163 ( L126gat_wire, L466gat, L517gat );
    nor2 U253 ( L341gat, L659gat, L731gat );
    nor2 U348 ( L334gat, L836gat, L845gat );
    and2 U274 ( L237gat_wire, L705gat, L752gat );
    nor2 U181 ( L318gat, L508gat, L539gat );
    nand2 U186 ( L518gat, L519gat, L544gat );
    nor2 U291 ( L736gat, L737gat, L769gat );
    nor2 U301 ( L757gat, L758gat, L786gat );
    nand3 U326 ( L741gat, L764gat, L813gat, L819gat );
    nor2 U296 ( L748gat, L749gat, L777gat );
    and2 U306 ( L708gat, L778gat, L791gat );
    nand4 U321 ( L805gat, L787gat, L731gat, L529gat, L811gat );
    buffer U368 ( L857gat, L865gat_wire );
    nand2 U38 ( L171gat_wire, L177gat_wire, L326gat );
    nor2 U143 ( L416gat, L445gat, L495gat );
    and2 U273 ( L228gat_wire, L708gat, L751gat );
    and2 U158 ( L146gat_wire, L483gat, L512gat );
    nand2 U164 ( L130gat_wire, L492gat, L518gat );
    nand2 U254 ( L654gat, L261gat_wire, L732gat );
    and2 U268 ( L237gat_wire, L687gat, L746gat );
    and2 U44 ( L210gat_wire, L91gat_wire, L332gat );
    or2 U56 ( L270gat, L273gat, L344gat );
    inv U94 ( L366gat, L408gat );
    and2 U136 ( L310gat, L432gat, L482gat );
    and2 U354 ( L219gat_wire, L842gat, L851gat );
    inv U373 ( L862gat, L870gat );
    and2 U206 ( L246gat_wire, L553gat, L596gat );
    nand2 U71 ( L305gat, L306gat, L363gat );
    and2 U221 ( L246gat_wire, L573gat, L640gat );
    and2 U111 ( L404gat, L405gat, L425gat );
    buffer U124 ( L403gat, L450gat_wire );
    or2 U214 ( L565gat, L177gat_wire, L619gat );
    inv U63 ( L293gat, L351gat );
    inv U233 ( L597gat, L670gat );
    and2 U86 ( L348gat, L73gat_wire, L400gat );
    and2 U103 ( L210gat_wire, L369gat, L417gat );
    inv U188 ( L530gat, L550gat );
    nor2 U328 ( L806gat, L807gat, L825gat );
    nor2 U346 ( L832gat, L833gat, L843gat );
    inv U361 ( L849gat, L858gat );
    and3 U16 ( L59gat_wire, L36gat_wire, L80gat_wire, L295gat );
    and2 U31 ( L17gat_wire, L138gat_wire, L317gat );
    nor2 U151 ( L477gat, L478gat, L505gat );
    and2 U261 ( L228gat_wire, L673gat, L739gat );
    nand2 U176 ( L498gat, L499gat, L530gat );
    nand2 U78 ( L330gat, L331gat, L385gat );
    and2 U118 ( L411gat, L412gat, L444gat );
    nand2 U193 ( L538gat, L507gat, L561gat );
    and2 U246 ( L635gat, L632gat, L708gat );
    nand2 U284 ( L635gat, L713gat, L762gat );
    nor2 U333 ( L665gat, L815gat, L830gat );
    nor2 U314 ( L792gat, L793gat, L804gat );
    nor2 U228 ( L552gat, L588gat, L660gat );
endmodule

