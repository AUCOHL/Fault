module c3540(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,
  G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G3519,G3520,G3521,G3522,
  G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,
  G3535,G3536,G3537,G3538,G3539,G3540,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,
  G45,G46,G47,G48,G49,G5,G50,G6,G7,G8,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50;
output G3519,G3520,G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,
  G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540;

  wire G353,G363,G368,G377,G381,G384,G388,G397,G400,G404,G413,G422,G425,G434,
    G438,G447,G451,G461,G466,G467,G470,G477,G480,G484,G491,G492,G496,G501,G518,
    G519,G523,G527,G530,G533,G534,G537,G540,G543,G546,G549,G552,G556,G559,G562,
    G565,G568,G572,G575,G578,G581,G584,G587,G588,G589,G590,G593,G594,G611,G612,
    G613,G614,G615,G618,G621,G624,G627,G630,G633,G636,G639,G642,G645,G648,G651,
    G654,G657,G660,G663,G666,G667,G684,G685,G686,G691,G708,G713,G714,G715,G716,
    G717,G718,G719,G720,G721,G722,G723,G724,G725,G726,G727,G730,G731,G734,G735,
    G736,G739,G742,G745,G749,G753,G762,G769,G772,G775,G778,G781,G784,G785,G786,
    G787,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,G805,G810,G813,
    G816,G831,G848,G849,G850,G851,G852,G853,G854,G855,G856,G873,G874,G875,G882,
    G883,G884,G887,G890,G891,G892,G893,G894,G897,G898,G901,G904,G907,G910,G913,
    G916,G919,G922,G925,G928,G929,G930,G931,G932,G933,G934,G935,G939,G956,G957,
    G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,
    G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,G986,G989,
    G992,G993,G994,G995,G996,G997,G998,G999,G1000,G1001,G1002,G1003,G1004,
    G1005,G1008,G1011,G1012,G1015,G1016,G1017,G1018,G1019,G1020,G1021,G1022,
    G1023,G1024,G1025,G1034,G1043,G1048,G1051,G1052,G1053,G1054,G1055,G1056,
    G1057,G1058,G1059,G1060,G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,
    G1069,G1070,G1071,G1072,G1073,G1074,G1077,G1080,G1083,G1086,G1089,G1092,
    G1095,G1104,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,G1121,G1122,
    G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,
    G1135,G1136,G1137,G1140,G1141,G1142,G1145,G1146,G1147,G1150,G1151,G1152,
    G1155,G1156,G1157,G1160,G1161,G1162,G1165,G1166,G1167,G1170,G1171,G1172,
    G1175,G1176,G1179,G1180,G1184,G1189,G1193,G1197,G1200,G1203,G1206,G1207,
    G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,
    G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,
    G1234,G1235,G1236,G1237,G1238,G1239,G1240,G1241,G1242,G1243,G1244,G1249,
    G1258,G1263,G1272,G1275,G1278,G1281,G1284,G1287,G1290,G1293,G1296,G1297,
    G1298,G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,
    G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,
    G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1345,G1348,G1349,G1350,G1351,
    G1352,G1353,G1354,G1357,G1360,G1363,G1366,G1369,G1372,G1375,G1378,G1379,
    G1380,G1381,G1390,G1399,G1400,G1401,G1402,G1403,G1404,G1405,G1406,G1407,
    G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1418,G1421,G1424,G1427,
    G1430,G1433,G1436,G1439,G1442,G1445,G1448,G1451,G1454,G1457,G1460,G1463,
    G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,
    G1478,G1479,G1482,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,
    G1494,G1495,G1496,G1497,G1498,G1499,G1500,G1501,G1502,G1503,G1504,G1505,
    G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1517,G1518,G1519,
    G1520,G1521,G1522,G1523,G1524,G1527,G1528,G1529,G1538,G1547,G1556,G1565,
    G1574,G1583,G1592,G1601,G1610,G1619,G1628,G1637,G1646,G1655,G1664,G1673,
    G1674,G1675,G1676,G1677,G1678,G1679,G1680,G1681,G1682,G1683,G1684,G1685,
    G1686,G1687,G1688,G1689,G1693,G1697,G1700,G1703,G1707,G1711,G1714,G1718,
    G1722,G1725,G1729,G1733,G1738,G1743,G1747,G1751,G1756,G1760,G1764,G1769,
    G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,G1781,
    G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,
    G1794,G1795,G1796,G1799,G1802,G1805,G1806,G1807,G1808,G1809,G1810,G1811,
    G1812,G1813,G1816,G1819,G1823,G1826,G1827,G1828,G1829,G1830,G1831,G1832,
    G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,G1841,G1842,G1843,G1844,
    G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,
    G1857,G1858,G1859,G1860,G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,
    G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
    G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,
    G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,G1901,G1902,G1903,G1904,
    G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,
    G1917,G1918,G1919,G1920,G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,
    G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
    G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,
    G1953,G1954,G1955,G1958,G1961,G1962,G1965,G1968,G1971,G1974,G1977,G1978,
    G1981,G1984,G1985,G1988,G1991,G1992,G1995,G1998,G2001,G2004,G2007,G2008,
    G2011,G2014,G2015,G2018,G2021,G2024,G2027,G2030,G2033,G2034,G2035,G2036,
    G2037,G2038,G2039,G2040,G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,
    G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
    G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,
    G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,G2081,G2082,G2083,G2084,
    G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,
    G2097,G2098,G2099,G2100,G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,
    G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
    G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,
    G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,G2141,G2142,G2143,G2144,
    G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,
    G2157,G2158,G2159,G2160,G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,
    G2169,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,G2181,G2182,
    G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2195,G2198,
    G2199,G2200,G2204,G2208,G2211,G2214,G2215,G2216,G2219,G2222,G2223,G2224,
    G2227,G2230,G2231,G2232,G2236,G2240,G2243,G2246,G2247,G2248,G2251,G2254,
    G2255,G2256,G2257,G2260,G2263,G2266,G2269,G2272,G2275,G2278,G2281,G2284,
    G2287,G2290,G2293,G2296,G2299,G2302,G2305,G2308,G2311,G2312,G2313,G2314,
    G2315,G2316,G2317,G2318,G2319,G2320,G2321,G2322,G2323,G2324,G2325,G2326,
    G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,
    G2339,G2340,G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,
    G2351,G2352,G2353,G2354,G2355,G2356,G2359,G2362,G2363,G2364,G2365,G2368,
    G2369,G2372,G2373,G2374,G2375,G2378,G2381,G2382,G2383,G2384,G2387,G2388,
    G2391,G2392,G2393,G2396,G2397,G2398,G2399,G2400,G2401,G2404,G2405,G2406,
    G2407,G2408,G2411,G2414,G2415,G2416,G2417,G2418,G2419,G2420,G2421,G2422,
    G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2436,G2437,G2441,G2444,
    G2450,G2451,G2455,G2458,G2459,G2460,G2461,G2462,G2463,G2464,G2465,G2466,
    G2467,G2468,G2471,G2472,G2475,G2476,G2479,G2482,G2485,G2488,G2491,G2494,
    G2497,G2500,G2501,G2502,G2507,G2512,G2515,G2518,G2521,G2524,G2527,G2530,
    G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2542,G2543,G2546,
    G2547,G2550,G2551,G2552,G2556,G2557,G2558,G2561,G2562,G2563,G2566,G2569,
    G2570,G2571,G2574,G2577,G2580,G2583,G2586,G2589,G2592,G2595,G2598,G2601,
    G2604,G2607,G2610,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,G2623,
    G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,
    G2636,G2637,G2638,G2639,G2640,G2643,G2646,G2647,G2648,G2651,G2654,G2655,
    G2656,G2657,G2658,G2659,G2660,G2661,G2662,G2663,G2664,G2665,G2666,G2669,
    G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,G2681,G2682,G2683,G2684,
    G2685,G2686,G2687,G2690,G2693,G2694,G2697,G2698,G2699,G2705,G2708,G2711,
    G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,G2721,G2728,G2733,
    G2736,G2739,G2740,G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2750,G2753,
    G2759,G2763,G2768,G2773,G2778,G2779,G2780,G2781,G2784,G2787,G2788,G2789,
    G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2799,G2803,G2804,G2805,G2808,
    G2809,G2810,G2811,G2816,G2820,G2821,G2822,G2823,G2826,G2827,G2828,G2829,
    G2830,G2831,G2832,G2833,G2836,G2839,G2842,G2845,G2848,G2851,G2854,G2857,
    G2860,G2863,G2866,G2869,G2872,G2875,G2876,G2877,G2880,G2883,G2884,G2887,
    G2890,G2893,G2896,G2899,G2902,G2905,G2906,G2909,G2910,G2911,G2912,G2913,
    G2916,G2917,G2918,G2919,G2920,G2923,G2926,G2929,G2932,G2935,G2936,G2937,
    G2938,G2939,G2942,G2943,G2944,G2947,G2950,G2951,G2952,G2953,G2954,G2955,
    G2956,G2957,G2958,G2959,G2960,G2961,G2962,G2965,G2968,G2971,G2974,G2975,
    G2978,G2979,G2980,G2981,G2984,G2985,G2986,G2990,G2991,G2994,G2995,G2996,
    G2999,G3002,G3005,G3006,G3007,G3010,G3011,G3012,G3015,G3016,G3017,G3018,
    G3021,G3024,G3027,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,
    G3039,G3042,G3045,G3048,G3051,G3054,G3057,G3058,G3059,G3060,G3061,G3062,
    G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3072,G3075,G3078,G3081,G3082,
    G3083,G3084,G3085,G3086,G3089,G3090,G3094,G3095,G3099,G3100,G3103,G3106,
    G3107,G3110,G3114,G3115,G3116,G3117,G3118,G3119,G3120,G3121,G3122,G3126,
    G3129,G3132,G3135,G3136,G3137,G3138,G3139,G3140,G3143,G3146,G3149,G3152,
    G3155,G3158,G3159,G3160,G3164,G3165,G3168,G3169,G3170,G3171,G3174,G3177,
    G3180,G3183,G3186,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3199,G3202,
    G3203,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,
    G3217,G3220,G3223,G3226,G3227,G3230,G3231,G3232,G3233,G3234,G3235,G3236,
    G3237,G3240,G3243,G3246,G3247,G3248,G3249,G3250,G3251,G3254,G3257,G3258,
    G3259,G3260,G3261,G3262,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,
    G3275,G3278,G3281,G3284,G3287,G3288,G3291,G3294,G3297,G3300,G3301,G3302,
    G3305,G3308,G3311,G3312,G3317,G3320,G3323,G3326,G3329,G3332,G3337,G3340,
    G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3350,G3353,G3356,G3359,G3360,
    G3363,G3366,G3367,G3370,G3373,G3376,G3379,G3380,G3383,G3386,G3387,G3388,
    G3391,G3394,G3395,G3396,G3399,G3402,G3403,G3404,G3405,G3406,G3407,G3408,
    G3409,G3412,G3415,G3416,G3417,G3418,G3419,G3420,G3421,G3422,G3423,G3424,
    G3425,G3428,G3429,G3430,G3431,G3432,G3436,G3437,G3438,G3439,G3440,G3441,
    G3444,G3445,G3448,G3449,G3452,G3453,G3456,G3459,G3460,G3461,G3464,G3465,
    G3466,G3467,G3468,G3471,G3474,G3475,G3478,G3481,G3484,G3487,G3488,G3489,
    G3490,G3491,G3494,G3497,G3500,G3503,G3504,G3505,G3506,G3507,G3508,G3509,
    G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518;

  not NOT_0(G353,G7);
  not NOT_1(G363,G7);
  not NOT_2(G368,G8);
  not NOT_3(G377,G8);
  not NOT_4(G381,G9);
  not NOT_5(G384,G9);
  not NOT_6(G388,G9);
  not NOT_7(G397,G10);
  not NOT_8(G400,G10);
  not NOT_9(G404,G10);
  not NOT_10(G413,G11);
  not NOT_11(G422,G11);
  not NOT_12(G425,G12);
  not NOT_13(G434,G12);
  not NOT_14(G438,G13);
  not NOT_15(G447,G13);
  not NOT_16(G451,G14);
  not NOT_17(G461,G14);
  or OR2_0(G466,G35,G36);
  not NOT_18(G467,G1);
  not NOT_19(G470,G1);
  not NOT_20(G477,G1);
  not NOT_21(G480,G2);
  not NOT_22(G484,G2);
  and AND2_0(G491,G2,G3);
  not NOT_23(G492,G3);
  not NOT_24(G496,G3);
  not NOT_25(G501,G3);
  not NOT_26(G518,G4);
  not NOT_27(G519,G4);
  not NOT_28(G523,G4);
  and AND2_1(G527,G4,G5);
  not NOT_29(G530,G5);
  or OR2_1(G533,G5,G6);
  not NOT_30(G534,G6);
  not NOT_31(G537,G6);
  not NOT_32(G540,G7);
  not NOT_33(G543,G8);
  not NOT_34(G546,G8);
  not NOT_35(G549,G9);
  not NOT_36(G552,G9);
  not NOT_37(G556,G11);
  not NOT_38(G559,G11);
  not NOT_39(G562,G12);
  not NOT_40(G565,G12);
  not NOT_41(G568,G13);
  not NOT_42(G572,G1);
  not NOT_43(G575,G9);
  not NOT_44(G578,G13);
  not NOT_45(G581,G3);
  not NOT_46(G584,G25);
  not NOT_47(G587,G26);
  and AND2_2(G588,G3,G26);
  nand NAND2_0(G589,G3,G26);
  and AND2_3(G590,G3,G24);
  not NOT_48(G593,G3);
  or OR2_2(G594,G49,G4);
  nand NAND2_1(G611,G1,G2);
  nand NAND3_0(G612,G1,G3,G4);
  not NOT_49(G613,G3);
  not NOT_50(G614,G4);
  not NOT_51(G615,G24);
  not NOT_52(G618,G27);
  not NOT_53(G621,G48);
  not NOT_54(G624,G30);
  not NOT_55(G627,G31);
  not NOT_56(G630,G32);
  not NOT_57(G633,G33);
  not NOT_58(G636,G34);
  not NOT_59(G639,G35);
  not NOT_60(G642,G36);
  not NOT_61(G645,G37);
  not NOT_62(G648,G7);
  not NOT_63(G651,G8);
  not NOT_64(G654,G8);
  not NOT_65(G657,G12);
  not NOT_66(G660,G12);
  not NOT_67(G663,G47);
  and AND2_4(G666,G34,G466);
  or OR2_3(G667,G518,G3);
  or OR2_4(G684,G593,G23);
  not NOT_68(G685,G491);
  or OR2_5(G686,G613,G1);
  and AND2_5(G691,G611,G612);
  or OR2_6(G708,G614,G1);
  and AND3_0(G713,G540,G546,G552);
  nand NAND2_2(G714,G30,G353);
  nand NAND2_3(G715,G31,G368);
  nand NAND2_4(G716,G32,G388);
  nand NAND2_5(G717,G33,G404);
  nand NAND2_6(G718,G34,G413);
  nand NAND2_7(G719,G35,G425);
  nand NAND2_8(G720,G36,G438);
  nand NAND2_9(G721,G37,G451);
  not NOT_69(G722,G624);
  not NOT_70(G723,G627);
  not NOT_71(G724,G630);
  not NOT_72(G725,G633);
  nand NAND2_10(G726,G377,G384);
  nand NAND2_11(G727,G434,G447);
  nand NAND2_12(G730,G381,G397);
  not NOT_73(G731,G363);
  not NOT_74(G734,G651);
  not NOT_75(G735,G657);
  not NOT_76(G736,G537);
  not NOT_77(G739,G537);
  not NOT_78(G742,G480);
  not NOT_79(G745,G523);
  not NOT_80(G749,G530);
  and AND2_6(G753,G477,G533);
  and AND3_1(G762,G477,G534,G530);
  and AND2_7(G769,G467,G534);
  and AND3_2(G772,G470,G484,G496);
  nand NAND3_1(G775,G470,G484,G496);
  nand NAND2_13(G778,G470,G484);
  not NOT_81(G781,G572);
  nand NAND3_2(G784,G480,G492,G6);
  nand NAND3_3(G785,G540,G546,G552);
  not NOT_82(G786,G654);
  and AND3_3(G787,G559,G565,G568);
  nand NAND3_4(G790,G559,G565,G568);
  not NOT_83(G791,G660);
  not NOT_84(G792,G501);
  not NOT_85(G793,G501);
  not NOT_86(G794,G501);
  not NOT_87(G795,G501);
  not NOT_88(G796,G501);
  not NOT_89(G797,G501);
  not NOT_90(G798,G501);
  not NOT_91(G799,G501);
  or OR2_7(G800,G581,G584);
  nor NOR2_0(G805,G581,G584);
  not NOT_92(G810,G590);
  not NOT_93(G813,G590);
  not NOT_94(G816,G519);
  not NOT_95(G831,G523);
  not NOT_96(G848,G594);
  not NOT_97(G849,G594);
  not NOT_98(G850,G594);
  not NOT_99(G851,G594);
  not NOT_100(G852,G594);
  not NOT_101(G853,G594);
  not NOT_102(G854,G594);
  not NOT_103(G855,G594);
  or OR2_8(G856,G1,G685);
  not NOT_104(G873,G527);
  not NOT_105(G874,G527);
  and AND3_4(G875,G467,G480,G492);
  not NOT_106(G882,G615);
  not NOT_107(G883,G663);
  or OR2_9(G884,G618,G621);
  nor NOR2_1(G887,G618,G621);
  not NOT_108(G890,G636);
  not NOT_109(G891,G639);
  not NOT_110(G892,G642);
  not NOT_111(G893,G645);
  not NOT_112(G894,G377);
  not NOT_113(G897,G648);
  not NOT_114(G898,G384);
  not NOT_115(G901,G400);
  not NOT_116(G904,G422);
  not NOT_117(G907,G434);
  not NOT_118(G910,G447);
  not NOT_119(G913,G461);
  not NOT_120(G916,G575);
  not NOT_121(G919,G575);
  not NOT_122(G922,G578);
  not NOT_123(G925,G578);
  nand NAND2_14(G928,G400,G713);
  and AND4_0(G929,G714,G715,G716,G717);
  and AND4_1(G930,G718,G719,G720,G721);
  nand NAND2_15(G931,G627,G722);
  nand NAND2_16(G932,G624,G723);
  nand NAND2_17(G933,G633,G724);
  nand NAND2_18(G934,G630,G725);
  and AND2_8(G935,G353,G726);
  and AND2_9(G939,G572,G784);
  not NOT_124(G956,G667);
  and AND2_10(G957,G501,G667);
  and AND2_11(G958,G785,G792);
  not NOT_125(G959,G667);
  and AND2_12(G960,G501,G667);
  not NOT_126(G961,G667);
  and AND2_13(G962,G501,G667);
  and AND2_14(G963,G552,G794);
  not NOT_127(G964,G667);
  and AND2_15(G965,G501,G667);
  and AND2_16(G966,G10,G795);
  not NOT_128(G967,G667);
  and AND2_17(G968,G501,G667);
  and AND2_18(G969,G790,G796);
  not NOT_129(G970,G667);
  and AND2_19(G971,G501,G667);
  not NOT_130(G972,G667);
  and AND2_20(G973,G501,G667);
  and AND2_21(G974,G568,G798);
  not NOT_131(G975,G667);
  and AND2_22(G976,G501,G667);
  and AND2_23(G977,G14,G799);
  and AND2_24(G978,G28,G848);
  and AND2_25(G979,G29,G849);
  and AND2_26(G980,G30,G850);
  and AND2_27(G981,G31,G851);
  and AND2_28(G982,G32,G852);
  and AND2_29(G983,G33,G853);
  and AND2_30(G984,G34,G854);
  and AND2_31(G985,G35,G855);
  and AND3_5(G986,G1,G2,G873);
  and AND3_6(G989,G1,G2,G874);
  not NOT_132(G992,G691);
  not NOT_133(G993,G691);
  not NOT_134(G994,G691);
  not NOT_135(G995,G691);
  not NOT_136(G996,G691);
  not NOT_137(G997,G691);
  not NOT_138(G998,G691);
  not NOT_139(G999,G691);
  nand NAND2_19(G1000,G639,G890);
  nand NAND2_20(G1001,G636,G891);
  nand NAND2_21(G1002,G645,G892);
  nand NAND2_22(G1003,G642,G893);
  and AND2_32(G1004,G11,G727);
  nand NAND2_23(G1005,G931,G932);
  nand NAND2_24(G1008,G933,G934);
  nand NAND2_25(G1011,G929,G930);
  and AND2_33(G1012,G461,G787);
  nand NAND2_26(G1015,G461,G787);
  not NOT_140(G1016,G731);
  nand NAND2_27(G1017,G916,G734);
  not NOT_141(G1018,G916);
  and AND2_34(G1019,G381,G731);
  nand NAND2_28(G1020,G922,G735);
  not NOT_142(G1021,G922);
  nand NAND2_29(G1022,G11,G727);
  not NOT_143(G1023,G736);
  not NOT_144(G1024,G739);
  nand NAND2_30(G1025,G772,G519);
  nand NAND2_31(G1034,G772,G523);
  nand NAND3_5(G1043,G470,G742,G496);
  nand NAND4_0(G1048,G470,G484,G496,G749);
  nand NAND2_32(G1051,G919,G786);
  not NOT_145(G1052,G919);
  nand NAND2_33(G1053,G925,G791);
  not NOT_146(G1054,G925);
  not NOT_147(G1055,G775);
  not NOT_148(G1056,G781);
  not NOT_149(G1057,G778);
  and AND2_35(G1058,G543,G956);
  and AND2_36(G1059,G21,G957);
  and AND2_37(G1060,G549,G959);
  and AND2_38(G1061,G22,G960);
  and AND2_39(G1062,G10,G961);
  and AND2_40(G1063,G7,G962);
  and AND2_41(G1064,G556,G964);
  and AND2_42(G1065,G543,G965);
  and AND2_43(G1066,G562,G967);
  and AND2_44(G1067,G549,G968);
  and AND2_45(G1068,G13,G970);
  and AND2_46(G1069,G10,G971);
  and AND2_47(G1070,G14,G972);
  and AND2_48(G1071,G556,G973);
  and AND2_49(G1072,G39,G975);
  and AND2_50(G1073,G562,G976);
  and AND2_51(G1074,G26,G810);
  and AND2_52(G1077,G587,G810);
  and AND2_53(G1080,G588,G813);
  and AND2_54(G1083,G589,G813);
  nand NAND2_34(G1086,G745,G749);
  nand NAND2_35(G1089,G519,G749);
  nand NAND3_6(G1092,G470,G742,G684);
  nand NAND3_7(G1095,G484,G492,G745);
  nand NAND2_36(G1104,G484,G745);
  not NOT_150(G1113,G816);
  not NOT_151(G1114,G816);
  not NOT_152(G1115,G816);
  not NOT_153(G1116,G816);
  not NOT_154(G1117,G816);
  not NOT_155(G1118,G816);
  not NOT_156(G1119,G816);
  not NOT_157(G1120,G831);
  and AND2_55(G1121,G831,G594);
  not NOT_158(G1122,G831);
  and AND2_56(G1123,G831,G594);
  not NOT_159(G1124,G831);
  and AND2_57(G1125,G831,G594);
  not NOT_160(G1126,G831);
  and AND2_58(G1127,G831,G594);
  not NOT_161(G1128,G831);
  and AND2_59(G1129,G831,G594);
  not NOT_162(G1130,G831);
  and AND2_60(G1131,G831,G594);
  not NOT_163(G1132,G831);
  and AND2_61(G1133,G831,G594);
  not NOT_164(G1134,G831);
  and AND2_62(G1135,G831,G594);
  and AND2_63(G1136,G691,G856);
  nor NOR2_2(G1137,G7,G856);
  not NOT_165(G1140,G753);
  and AND2_64(G1141,G691,G856);
  nor NOR2_3(G1142,G8,G856);
  not NOT_166(G1145,G753);
  and AND2_65(G1146,G691,G856);
  nor NOR2_4(G1147,G9,G856);
  not NOT_167(G1150,G753);
  and AND2_66(G1151,G691,G856);
  nor NOR2_5(G1152,G10,G856);
  not NOT_168(G1155,G753);
  and AND2_67(G1156,G691,G856);
  nor NOR2_6(G1157,G11,G856);
  not NOT_169(G1160,G769);
  and AND2_68(G1161,G691,G856);
  nor NOR2_7(G1162,G12,G856);
  not NOT_170(G1165,G762);
  and AND2_69(G1166,G691,G856);
  nor NOR2_8(G1167,G13,G856);
  not NOT_171(G1170,G762);
  and AND2_70(G1171,G691,G856);
  nor NOR2_9(G1172,G14,G856);
  not NOT_172(G1175,G762);
  and AND2_71(G1176,G875,G27);
  nand NAND2_37(G1179,G875,G27);
  and AND3_7(G1180,G875,G27,G48);
  nand NAND3_8(G1184,G875,G27,G48);
  and AND3_8(G1189,G875,G27,G48);
  nand NAND3_9(G1193,G875,G27,G48);
  not NOT_173(G1197,G887);
  nand NAND2_38(G1200,G1000,G1001);
  nand NAND2_39(G1203,G1002,G1003);
  not NOT_174(G1206,G894);
  nand NAND2_40(G1207,G894,G897);
  not NOT_175(G1208,G898);
  not NOT_176(G1209,G901);
  not NOT_177(G1210,G904);
  not NOT_178(G1211,G907);
  not NOT_179(G1212,G910);
  not NOT_180(G1213,G913);
  nand NAND2_41(G1214,G651,G1018);
  nand NAND2_42(G1215,G657,G1021);
  and AND2_72(G1216,G935,G739);
  nand NAND2_43(G1217,G654,G1052);
  nand NAND2_44(G1218,G660,G1054);
  and AND2_73(G1219,G666,G1055);
  or OR3_0(G1222,G958,G1058,G1059);
  or OR3_1(G1223,G963,G1062,G1063);
  or OR3_2(G1224,G966,G1064,G1065);
  or OR3_3(G1225,G969,G1066,G1067);
  or OR3_4(G1226,G974,G1070,G1071);
  or OR3_5(G1227,G977,G1072,G1073);
  and AND2_74(G1228,G10,G1120);
  and AND2_75(G1229,G29,G1121);
  and AND2_76(G1230,G11,G1122);
  and AND2_77(G1231,G30,G1123);
  and AND2_78(G1232,G12,G1124);
  and AND2_79(G1233,G31,G1125);
  and AND2_80(G1234,G13,G1126);
  and AND2_81(G1235,G32,G1127);
  and AND2_82(G1236,G14,G1128);
  and AND2_83(G1237,G33,G1129);
  and AND2_84(G1238,G39,G1130);
  and AND2_85(G1239,G34,G1131);
  and AND2_86(G1240,G40,G1132);
  and AND2_87(G1241,G35,G1133);
  and AND2_88(G1242,G41,G1134);
  and AND2_89(G1243,G36,G1135);
  not NOT_181(G1244,G986);
  not NOT_182(G1249,G986);
  not NOT_183(G1258,G989);
  not NOT_184(G1263,G989);
  and AND3_9(G1272,G7,G686,G1136);
  and AND3_10(G1275,G8,G686,G1141);
  and AND3_11(G1278,G9,G686,G1146);
  and AND3_12(G1281,G10,G686,G1151);
  and AND3_13(G1284,G11,G708,G1156);
  and AND3_14(G1287,G12,G708,G1161);
  and AND3_15(G1290,G13,G708,G1166);
  and AND3_16(G1293,G14,G708,G1171);
  not NOT_185(G1296,G939);
  not NOT_186(G1297,G939);
  not NOT_187(G1298,G939);
  not NOT_188(G1299,G939);
  not NOT_189(G1300,G939);
  not NOT_190(G1301,G939);
  not NOT_191(G1302,G939);
  not NOT_192(G1303,G939);
  nand NAND2_45(G1304,G648,G1206);
  nand NAND2_46(G1305,G901,G1208);
  nand NAND2_47(G1306,G898,G1209);
  nand NAND2_48(G1307,G907,G1210);
  nand NAND2_49(G1308,G904,G1211);
  nand NAND2_50(G1309,G913,G1212);
  nand NAND2_51(G1310,G910,G1213);
  not NOT_193(G1311,G1200);
  not NOT_194(G1312,G1203);
  not NOT_195(G1313,G1025);
  and AND2_90(G1314,G1025,G1034);
  not NOT_196(G1315,G1034);
  nand NAND2_52(G1316,G1017,G1214);
  nand NAND2_53(G1317,G1020,G1215);
  and AND4_2(G1318,G1012,G730,G363,G8);
  not NOT_197(G1319,G1025);
  and AND2_91(G1320,G1025,G1034);
  not NOT_198(G1321,G1034);
  not NOT_199(G1322,G1025);
  not NOT_200(G1323,G1034);
  and AND2_92(G1324,G1025,G1034);
  not NOT_201(G1325,G1025);
  not NOT_202(G1326,G1034);
  and AND2_93(G1327,G1025,G1034);
  not NOT_203(G1328,G1048);
  not NOT_204(G1345,G1048);
  nand NAND2_54(G1348,G1051,G1217);
  nand NAND2_55(G1349,G1053,G1218);
  not NOT_205(G1350,G1043);
  and AND2_94(G1351,G1043,G775);
  not NOT_206(G1352,G1043);
  and AND2_95(G1353,G778,G1043);
  nand NAND2_56(G1354,G805,G1083);
  nand NAND2_57(G1357,G805,G1080);
  nand NAND2_58(G1360,G800,G1083);
  nand NAND2_59(G1363,G800,G1080);
  nand NAND2_60(G1366,G805,G1077);
  nand NAND2_61(G1369,G805,G1074);
  nand NAND2_62(G1372,G800,G1077);
  nand NAND2_63(G1375,G800,G1074);
  not NOT_207(G1378,G1086);
  not NOT_208(G1379,G1089);
  and AND2_96(G1380,G1086,G1089);
  not NOT_209(G1381,G1092);
  not NOT_210(G1390,G1092);
  not NOT_211(G1399,G1104);
  not NOT_212(G1400,G1104);
  not NOT_213(G1401,G1104);
  not NOT_214(G1402,G1104);
  not NOT_215(G1403,G1095);
  not NOT_216(G1404,G1095);
  not NOT_217(G1405,G1095);
  not NOT_218(G1406,G1095);
  or OR3_6(G1407,G1228,G978,G1229);
  or OR3_7(G1408,G1230,G979,G1231);
  or OR3_8(G1409,G1232,G980,G1233);
  or OR3_9(G1410,G1234,G981,G1235);
  or OR3_10(G1411,G1236,G982,G1237);
  or OR3_11(G1412,G1238,G983,G1239);
  or OR3_12(G1413,G1240,G984,G1241);
  or OR3_13(G1414,G1242,G985,G1243);
  and AND2_97(G1415,G1222,G992);
  and AND2_98(G1418,G1223,G994);
  and AND2_99(G1421,G1224,G995);
  and AND2_100(G1424,G1225,G996);
  and AND2_101(G1427,G1226,G998);
  and AND2_102(G1430,G1227,G999);
  not NOT_219(G1433,G1184);
  and AND2_103(G1436,G1197,G50);
  nand NAND2_64(G1439,G1197,G50);
  not NOT_220(G1442,G1005);
  not NOT_221(G1445,G1008);
  not NOT_222(G1448,G1005);
  not NOT_223(G1451,G1008);
  nand NAND2_65(G1454,G1207,G1304);
  nand NAND2_66(G1457,G1305,G1306);
  nand NAND2_67(G1460,G1307,G1308);
  nand NAND2_68(G1463,G1309,G1310);
  nand NAND2_69(G1466,G1203,G1311);
  nand NAND2_70(G1467,G1200,G1312);
  and AND2_104(G1468,G422,G1314);
  and AND3_17(G1469,G1316,G397,G1016);
  and AND2_105(G1470,G451,G1317);
  and AND2_106(G1471,G1318,G736);
  and AND2_107(G1472,G434,G1320);
  and AND2_108(G1473,G1022,G1323);
  and AND2_109(G1474,G461,G1324);
  and AND2_110(G1475,G1015,G1326);
  and AND2_111(G1476,G447,G1327);
  not NOT_224(G1477,G1348);
  not NOT_225(G1478,G1349);
  and AND2_112(G1479,G935,G1350);
  and AND2_113(G1482,G1011,G1351);
  and AND2_114(G1485,G363,G1380);
  and AND3_18(G1486,G1263,G30,G1140);
  and AND3_19(G1487,G1263,G38,G753);
  and AND2_115(G1488,G1258,G1407);
  and AND3_20(G1489,G1263,G31,G1145);
  and AND3_21(G1490,G1263,G38,G753);
  and AND2_116(G1491,G1258,G1408);
  and AND3_22(G1492,G1263,G32,G1150);
  and AND3_23(G1493,G1263,G38,G753);
  and AND2_117(G1494,G1258,G1409);
  and AND3_24(G1495,G1263,G33,G1155);
  and AND3_25(G1496,G1263,G38,G753);
  and AND2_118(G1497,G1258,G1410);
  and AND3_26(G1498,G1249,G34,G1160);
  and AND3_27(G1499,G1249,G38,G769);
  and AND2_119(G1500,G1244,G1411);
  and AND3_28(G1501,G1249,G35,G1165);
  and AND3_29(G1502,G1249,G38,G762);
  and AND2_120(G1503,G1244,G1412);
  and AND3_30(G1504,G1249,G36,G1170);
  and AND3_31(G1505,G1249,G38,G762);
  and AND2_121(G1506,G1244,G1413);
  and AND3_32(G1507,G1249,G37,G1175);
  and AND3_33(G1508,G1249,G38,G762);
  and AND2_122(G1509,G1244,G1414);
  not NOT_226(G1510,G1442);
  not NOT_227(G1511,G1445);
  not NOT_228(G1512,G1448);
  not NOT_229(G1513,G1451);
  nand NAND2_71(G1514,G1466,G1467);
  not NOT_230(G1517,G1454);
  not NOT_231(G1518,G1457);
  not NOT_232(G1519,G1460);
  not NOT_233(G1520,G1463);
  or OR2_10(G1521,G1469,G1019);
  not NOT_234(G1522,G1345);
  and AND2_123(G1523,G1345,G781);
  and AND2_124(G1524,G1470,G1352);
  and AND2_125(G1527,G1477,G793);
  and AND2_126(G1528,G1478,G797);
  not NOT_235(G1529,G1354);
  not NOT_236(G1538,G1357);
  not NOT_237(G1547,G1360);
  not NOT_238(G1556,G1363);
  not NOT_239(G1565,G1366);
  not NOT_240(G1574,G1369);
  not NOT_241(G1583,G1372);
  not NOT_242(G1592,G1375);
  not NOT_243(G1601,G1354);
  not NOT_244(G1610,G1357);
  not NOT_245(G1619,G1360);
  not NOT_246(G1628,G1363);
  not NOT_247(G1637,G1366);
  not NOT_248(G1646,G1369);
  not NOT_249(G1655,G1372);
  not NOT_250(G1664,G1375);
  not NOT_251(G1673,G1381);
  and AND2_127(G1674,G1381,G1104);
  not NOT_252(G1675,G1381);
  and AND2_128(G1676,G1381,G1104);
  not NOT_253(G1677,G1381);
  and AND2_129(G1678,G1381,G1104);
  not NOT_254(G1679,G1381);
  and AND2_130(G1680,G1381,G1104);
  not NOT_255(G1681,G1390);
  and AND2_131(G1682,G1390,G1095);
  not NOT_256(G1683,G1390);
  and AND2_132(G1684,G1390,G1095);
  not NOT_257(G1685,G1390);
  and AND2_133(G1686,G1390,G1095);
  not NOT_258(G1687,G1390);
  and AND2_134(G1688,G1390,G1095);
  or OR3_14(G1689,G1415,G1137,G1272);
  nor NOR3_0(G1693,G1415,G1137,G1272);
  or OR3_15(G1697,G1486,G1487,G1488);
  or OR3_16(G1700,G1489,G1490,G1491);
  or OR3_17(G1703,G1418,G1147,G1278);
  nor NOR3_1(G1707,G1418,G1147,G1278);
  or OR3_18(G1711,G1492,G1493,G1494);
  or OR3_19(G1714,G1421,G1152,G1281);
  nor NOR3_2(G1718,G1421,G1152,G1281);
  or OR3_20(G1722,G1495,G1496,G1497);
  or OR3_21(G1725,G1424,G1157,G1284);
  nor NOR3_3(G1729,G1424,G1157,G1284);
  or OR3_22(G1733,G1498,G1499,G1500);
  or OR3_23(G1738,G1501,G1502,G1503);
  or OR3_24(G1743,G1427,G1167,G1290);
  nor NOR3_4(G1747,G1427,G1167,G1290);
  or OR3_25(G1751,G1504,G1505,G1506);
  or OR3_26(G1756,G1430,G1172,G1293);
  nor NOR3_5(G1760,G1430,G1172,G1293);
  or OR3_27(G1764,G1507,G1508,G1509);
  not NOT_259(G1769,G1433);
  not NOT_260(G1770,G1328);
  and AND2_135(G1771,G939,G1328);
  not NOT_261(G1772,G1328);
  and AND2_136(G1773,G939,G1328);
  not NOT_262(G1774,G1328);
  and AND2_137(G1775,G939,G1328);
  not NOT_263(G1776,G1328);
  and AND2_138(G1777,G939,G1328);
  not NOT_264(G1778,G1328);
  and AND2_139(G1779,G939,G1328);
  not NOT_265(G1780,G1328);
  and AND2_140(G1781,G939,G1328);
  not NOT_266(G1782,G1328);
  and AND2_141(G1783,G939,G1328);
  not NOT_267(G1784,G1328);
  and AND2_142(G1785,G939,G1328);
  or OR3_28(G1786,G1479,G1219,G1482);
  nor NOR3_6(G1787,G1479,G1219,G1482);
  nand NAND2_72(G1788,G1445,G1510);
  nand NAND2_73(G1789,G1442,G1511);
  nand NAND2_74(G1790,G1451,G1512);
  nand NAND2_75(G1791,G1448,G1513);
  nand NAND2_76(G1792,G1457,G1517);
  nand NAND2_77(G1793,G1454,G1518);
  nand NAND2_78(G1794,G1463,G1519);
  nand NAND2_79(G1795,G1460,G1520);
  and AND2_143(G1796,G935,G1522);
  and AND2_144(G1799,G1012,G1523);
  and AND2_145(G1802,G1521,G1057);
  or OR3_29(G1805,G1527,G1060,G1061);
  or OR3_30(G1806,G1528,G1068,G1069);
  and AND2_146(G1807,G363,G1674);
  and AND2_147(G1808,G377,G1676);
  and AND2_148(G1809,G384,G1678);
  and AND2_149(G1810,G400,G1680);
  not NOT_268(G1811,G1787);
  nand NAND2_80(G1812,G1788,G1789);
  nand NAND2_81(G1813,G1790,G1791);
  not NOT_269(G1816,G1514);
  nand NAND2_82(G1819,G1792,G1793);
  nand NAND2_83(G1823,G1794,G1795);
  and AND2_150(G1826,G1514,G1313);
  not NOT_270(G1827,G1529);
  not NOT_271(G1828,G1538);
  not NOT_272(G1829,G1547);
  not NOT_273(G1830,G1556);
  not NOT_274(G1831,G1565);
  not NOT_275(G1832,G1574);
  not NOT_276(G1833,G1583);
  not NOT_277(G1834,G1592);
  not NOT_278(G1835,G1529);
  not NOT_279(G1836,G1538);
  not NOT_280(G1837,G1547);
  not NOT_281(G1838,G1556);
  not NOT_282(G1839,G1565);
  not NOT_283(G1840,G1574);
  not NOT_284(G1841,G1583);
  not NOT_285(G1842,G1592);
  not NOT_286(G1843,G1529);
  not NOT_287(G1844,G1538);
  not NOT_288(G1845,G1547);
  not NOT_289(G1846,G1556);
  not NOT_290(G1847,G1565);
  not NOT_291(G1848,G1574);
  not NOT_292(G1849,G1583);
  not NOT_293(G1850,G1592);
  not NOT_294(G1851,G1529);
  not NOT_295(G1852,G1538);
  not NOT_296(G1853,G1547);
  not NOT_297(G1854,G1556);
  not NOT_298(G1855,G1565);
  not NOT_299(G1856,G1574);
  not NOT_300(G1857,G1583);
  not NOT_301(G1858,G1592);
  not NOT_302(G1859,G1529);
  not NOT_303(G1860,G1538);
  not NOT_304(G1861,G1547);
  not NOT_305(G1862,G1556);
  not NOT_306(G1863,G1565);
  not NOT_307(G1864,G1574);
  not NOT_308(G1865,G1583);
  not NOT_309(G1866,G1592);
  not NOT_310(G1867,G1529);
  not NOT_311(G1868,G1538);
  not NOT_312(G1869,G1547);
  not NOT_313(G1870,G1556);
  not NOT_314(G1871,G1565);
  not NOT_315(G1872,G1574);
  not NOT_316(G1873,G1583);
  not NOT_317(G1874,G1592);
  not NOT_318(G1875,G1529);
  not NOT_319(G1876,G1538);
  not NOT_320(G1877,G1547);
  not NOT_321(G1878,G1556);
  not NOT_322(G1879,G1565);
  not NOT_323(G1880,G1574);
  not NOT_324(G1881,G1583);
  not NOT_325(G1882,G1592);
  not NOT_326(G1883,G1529);
  not NOT_327(G1884,G1538);
  not NOT_328(G1885,G1547);
  not NOT_329(G1886,G1556);
  not NOT_330(G1887,G1565);
  not NOT_331(G1888,G1574);
  not NOT_332(G1889,G1583);
  not NOT_333(G1890,G1592);
  not NOT_334(G1891,G1601);
  not NOT_335(G1892,G1610);
  not NOT_336(G1893,G1619);
  not NOT_337(G1894,G1628);
  not NOT_338(G1895,G1637);
  not NOT_339(G1896,G1646);
  not NOT_340(G1897,G1655);
  not NOT_341(G1898,G1664);
  not NOT_342(G1899,G1601);
  not NOT_343(G1900,G1610);
  not NOT_344(G1901,G1619);
  not NOT_345(G1902,G1628);
  not NOT_346(G1903,G1637);
  not NOT_347(G1904,G1646);
  not NOT_348(G1905,G1655);
  not NOT_349(G1906,G1664);
  not NOT_350(G1907,G1601);
  not NOT_351(G1908,G1610);
  not NOT_352(G1909,G1619);
  not NOT_353(G1910,G1628);
  not NOT_354(G1911,G1637);
  not NOT_355(G1912,G1646);
  not NOT_356(G1913,G1655);
  not NOT_357(G1914,G1664);
  not NOT_358(G1915,G1601);
  not NOT_359(G1916,G1610);
  not NOT_360(G1917,G1619);
  not NOT_361(G1918,G1628);
  not NOT_362(G1919,G1637);
  not NOT_363(G1920,G1646);
  not NOT_364(G1921,G1655);
  not NOT_365(G1922,G1664);
  not NOT_366(G1923,G1601);
  not NOT_367(G1924,G1610);
  not NOT_368(G1925,G1619);
  not NOT_369(G1926,G1628);
  not NOT_370(G1927,G1637);
  not NOT_371(G1928,G1646);
  not NOT_372(G1929,G1655);
  not NOT_373(G1930,G1664);
  not NOT_374(G1931,G1601);
  not NOT_375(G1932,G1610);
  not NOT_376(G1933,G1619);
  not NOT_377(G1934,G1628);
  not NOT_378(G1935,G1637);
  not NOT_379(G1936,G1646);
  not NOT_380(G1937,G1655);
  not NOT_381(G1938,G1664);
  not NOT_382(G1939,G1601);
  not NOT_383(G1940,G1610);
  not NOT_384(G1941,G1619);
  not NOT_385(G1942,G1628);
  not NOT_386(G1943,G1637);
  not NOT_387(G1944,G1646);
  not NOT_388(G1945,G1655);
  not NOT_389(G1946,G1664);
  not NOT_390(G1947,G1601);
  not NOT_391(G1948,G1610);
  not NOT_392(G1949,G1619);
  not NOT_393(G1950,G1628);
  not NOT_394(G1951,G1637);
  not NOT_395(G1952,G1646);
  not NOT_396(G1953,G1655);
  not NOT_397(G1954,G1664);
  not NOT_398(G1955,G1697);
  not NOT_399(G1958,G1697);
  not NOT_400(G1961,G1693);
  and AND2_151(G1962,G1805,G993);
  not NOT_401(G1965,G1700);
  not NOT_402(G1968,G1700);
  not NOT_403(G1971,G1711);
  not NOT_404(G1974,G1711);
  not NOT_405(G1977,G1707);
  not NOT_406(G1978,G1722);
  not NOT_407(G1981,G1722);
  not NOT_408(G1984,G1718);
  not NOT_409(G1985,G1733);
  not NOT_410(G1988,G1733);
  not NOT_411(G1991,G1729);
  and AND2_152(G1992,G1806,G997);
  not NOT_412(G1995,G1738);
  not NOT_413(G1998,G1738);
  not NOT_414(G2001,G1751);
  not NOT_415(G2004,G1751);
  not NOT_416(G2007,G1747);
  not NOT_417(G2008,G1764);
  not NOT_418(G2011,G1764);
  not NOT_419(G2014,G1760);
  and AND2_153(G2015,G1176,G1689);
  and AND2_154(G2018,G1180,G1703);
  and AND2_155(G2021,G1180,G1714);
  and AND2_156(G2024,G1180,G1725);
  and AND2_157(G2027,G1189,G1743);
  and AND2_158(G2030,G1189,G1756);
  not NOT_420(G2033,G1733);
  not NOT_421(G2034,G1738);
  not NOT_422(G2035,G1751);
  not NOT_423(G2036,G1764);
  and AND5_0(G2037,G1733,G1738,G1751,G1764,G882);
  not NOT_424(G2038,G1812);
  or OR3_31(G2039,G1826,G1315,G1468);
  and AND2_159(G2040,G15,G1827);
  and AND2_160(G2041,G22,G1828);
  and AND2_161(G2042,G21,G1829);
  and AND2_162(G2043,G20,G1830);
  and AND2_163(G2044,G19,G1831);
  and AND2_164(G2045,G18,G1832);
  and AND2_165(G2046,G17,G1833);
  and AND2_166(G2047,G16,G1834);
  and AND2_167(G2048,G16,G1835);
  and AND2_168(G2049,G353,G1836);
  and AND2_169(G2050,G22,G1837);
  and AND2_170(G2051,G21,G1838);
  and AND2_171(G2052,G20,G1839);
  and AND2_172(G2053,G19,G1840);
  and AND2_173(G2054,G18,G1841);
  and AND2_174(G2055,G17,G1842);
  and AND2_175(G2056,G17,G1843);
  and AND2_176(G2057,G368,G1844);
  and AND2_177(G2058,G353,G1845);
  and AND2_178(G2059,G22,G1846);
  and AND2_179(G2060,G21,G1847);
  and AND2_180(G2061,G20,G1848);
  and AND2_181(G2062,G19,G1849);
  and AND2_182(G2063,G18,G1850);
  and AND2_183(G2064,G18,G1851);
  and AND2_184(G2065,G388,G1852);
  and AND2_185(G2066,G368,G1853);
  and AND2_186(G2067,G353,G1854);
  and AND2_187(G2068,G22,G1855);
  and AND2_188(G2069,G21,G1856);
  and AND2_189(G2070,G20,G1857);
  and AND2_190(G2071,G19,G1858);
  and AND2_191(G2072,G19,G1859);
  and AND2_192(G2073,G404,G1860);
  and AND2_193(G2074,G388,G1861);
  and AND2_194(G2075,G368,G1862);
  and AND2_195(G2076,G353,G1863);
  and AND2_196(G2077,G22,G1864);
  and AND2_197(G2078,G21,G1865);
  and AND2_198(G2079,G20,G1866);
  and AND2_199(G2080,G20,G1867);
  and AND2_200(G2081,G413,G1868);
  and AND2_201(G2082,G404,G1869);
  and AND2_202(G2083,G388,G1870);
  and AND2_203(G2084,G368,G1871);
  and AND2_204(G2085,G353,G1872);
  and AND2_205(G2086,G22,G1873);
  and AND2_206(G2087,G21,G1874);
  and AND2_207(G2088,G21,G1875);
  and AND2_208(G2089,G425,G1876);
  and AND2_209(G2090,G413,G1877);
  and AND2_210(G2091,G404,G1878);
  and AND2_211(G2092,G388,G1879);
  and AND2_212(G2093,G368,G1880);
  and AND2_213(G2094,G353,G1881);
  and AND2_214(G2095,G22,G1882);
  and AND2_215(G2096,G22,G1883);
  and AND2_216(G2097,G438,G1884);
  and AND2_217(G2098,G425,G1885);
  and AND2_218(G2099,G413,G1886);
  and AND2_219(G2100,G404,G1887);
  and AND2_220(G2101,G388,G1888);
  and AND2_221(G2102,G368,G1889);
  and AND2_222(G2103,G353,G1890);
  and AND2_223(G2104,G39,G1891);
  and AND2_224(G2105,G368,G1892);
  and AND2_225(G2106,G388,G1893);
  and AND2_226(G2107,G404,G1894);
  and AND2_227(G2108,G413,G1895);
  and AND2_228(G2109,G425,G1896);
  and AND2_229(G2110,G438,G1897);
  and AND2_230(G2111,G451,G1898);
  and AND2_231(G2112,G40,G1899);
  and AND2_232(G2113,G388,G1900);
  and AND2_233(G2114,G404,G1901);
  and AND2_234(G2115,G413,G1902);
  and AND2_235(G2116,G425,G1903);
  and AND2_236(G2117,G438,G1904);
  and AND2_237(G2118,G451,G1905);
  and AND2_238(G2119,G39,G1906);
  and AND2_239(G2120,G41,G1907);
  and AND2_240(G2121,G404,G1908);
  and AND2_241(G2122,G413,G1909);
  and AND2_242(G2123,G425,G1910);
  and AND2_243(G2124,G438,G1911);
  and AND2_244(G2125,G451,G1912);
  and AND2_245(G2126,G39,G1913);
  and AND2_246(G2127,G40,G1914);
  and AND2_247(G2128,G42,G1915);
  and AND2_248(G2129,G413,G1916);
  and AND2_249(G2130,G425,G1917);
  and AND2_250(G2131,G438,G1918);
  and AND2_251(G2132,G451,G1919);
  and AND2_252(G2133,G39,G1920);
  and AND2_253(G2134,G40,G1921);
  and AND2_254(G2135,G41,G1922);
  and AND2_255(G2136,G43,G1923);
  and AND2_256(G2137,G425,G1924);
  and AND2_257(G2138,G438,G1925);
  and AND2_258(G2139,G451,G1926);
  and AND2_259(G2140,G39,G1927);
  and AND2_260(G2141,G40,G1928);
  and AND2_261(G2142,G41,G1929);
  and AND2_262(G2143,G42,G1930);
  and AND2_263(G2144,G44,G1931);
  and AND2_264(G2145,G438,G1932);
  and AND2_265(G2146,G451,G1933);
  and AND2_266(G2147,G39,G1934);
  and AND2_267(G2148,G40,G1935);
  and AND2_268(G2149,G41,G1936);
  and AND2_269(G2150,G42,G1937);
  and AND2_270(G2151,G43,G1938);
  and AND2_271(G2152,G45,G1939);
  and AND2_272(G2153,G451,G1940);
  and AND2_273(G2154,G39,G1941);
  and AND2_274(G2155,G40,G1942);
  and AND2_275(G2156,G41,G1943);
  and AND2_276(G2157,G42,G1944);
  and AND2_277(G2158,G43,G1945);
  and AND2_278(G2159,G44,G1946);
  and AND2_279(G2160,G46,G1947);
  and AND2_280(G2161,G39,G1948);
  and AND2_281(G2162,G40,G1949);
  and AND2_282(G2163,G41,G1950);
  and AND2_283(G2164,G42,G1951);
  and AND2_284(G2165,G43,G1952);
  and AND2_285(G2166,G44,G1953);
  and AND2_286(G2167,G45,G1954);
  and AND5_1(G2168,G2033,G2034,G2035,G2036,G615);
  not NOT_425(G2169,G1823);
  and AND2_287(G2172,G2038,G1023);
  and AND2_288(G2173,G1823,G1319);
  and AND2_289(G2174,G1819,G1024);
  nor NOR8_0(G2175,G2040,G2041,G2042,G2043,G2044,G2045,G2046,G2047);
  nor NOR8_1(G2176,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055);
  nor NOR8_2(G2177,G2056,G2057,G2058,G2059,G2060,G2061,G2062,G2063);
  nor NOR8_3(G2178,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071);
  nor NOR8_4(G2179,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079);
  nor NOR8_5(G2180,G2080,G2081,G2082,G2083,G2084,G2085,G2086,G2087);
  nor NOR8_6(G2181,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095);
  nor NOR8_7(G2182,G2096,G2097,G2098,G2099,G2100,G2101,G2102,G2103);
  nor NOR8_8(G2183,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111);
  nor NOR8_9(G2184,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119);
  nor NOR8_10(G2185,G2120,G2121,G2122,G2123,G2124,G2125,G2126,G2127);
  nor NOR8_11(G2186,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135);
  nor NOR8_12(G2187,G2136,G2137,G2138,G2139,G2140,G2141,G2142,G2143);
  nor NOR8_13(G2188,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151);
  nor NOR8_14(G2189,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159);
  nor NOR8_15(G2190,G2160,G2161,G2162,G2163,G2164,G2165,G2166,G2167);
  and AND2_290(G2191,G2039,G1682);
  and AND3_34(G2192,G23,G1689,G1955);
  and AND3_35(G2195,G24,G1689,G1958);
  and AND3_36(G2198,G25,G1693,G1958);
  and AND3_37(G2199,G26,G1693,G1955);
  or OR3_32(G2200,G1962,G1142,G1275);
  nor NOR3_7(G2204,G1962,G1142,G1275);
  and AND3_38(G2208,G23,G1703,G1971);
  and AND3_39(G2211,G24,G1703,G1974);
  and AND3_40(G2214,G25,G1707,G1974);
  and AND3_41(G2215,G26,G1707,G1971);
  and AND3_42(G2216,G23,G1714,G1978);
  and AND3_43(G2219,G24,G1714,G1981);
  and AND3_44(G2222,G25,G1718,G1981);
  and AND3_45(G2223,G26,G1718,G1978);
  and AND3_46(G2224,G23,G1725,G1985);
  and AND3_47(G2227,G24,G1725,G1988);
  and AND3_48(G2230,G25,G1729,G1988);
  and AND3_49(G2231,G26,G1729,G1985);
  or OR3_33(G2232,G1992,G1162,G1287);
  nor NOR3_8(G2236,G1992,G1162,G1287);
  and AND3_50(G2240,G23,G1743,G2001);
  and AND3_51(G2243,G24,G1743,G2004);
  and AND3_52(G2246,G25,G1747,G2004);
  and AND3_53(G2247,G26,G1747,G2001);
  and AND3_54(G2248,G23,G1756,G2008);
  and AND3_55(G2251,G24,G1756,G2011);
  and AND3_56(G2254,G25,G1760,G2011);
  and AND3_57(G2255,G26,G1760,G2008);
  or OR2_11(G2256,G2037,G2168);
  not NOT_426(G2257,G1813);
  not NOT_427(G2260,G1816);
  not NOT_428(G2263,G1813);
  not NOT_429(G2266,G1816);
  not NOT_430(G2269,G1819);
  not NOT_431(G2272,G1819);
  not NOT_432(G2275,G2015);
  not NOT_433(G2278,G2015);
  not NOT_434(G2281,G2018);
  not NOT_435(G2284,G2018);
  not NOT_436(G2287,G2021);
  not NOT_437(G2290,G2021);
  not NOT_438(G2293,G2024);
  not NOT_439(G2296,G2024);
  not NOT_440(G2299,G2027);
  not NOT_441(G2302,G2027);
  not NOT_442(G2305,G2030);
  not NOT_443(G2308,G2030);
  nor NOR2_10(G2311,G2172,G1471);
  or OR3_34(G2312,G2173,G1321,G1472);
  nor NOR2_11(G2313,G2174,G1216);
  and AND2_291(G2314,G2175,G1378);
  and AND2_292(G2315,G2183,G1379);
  and AND2_293(G2316,G2176,G1113);
  and AND2_294(G2317,G2184,G816);
  and AND2_295(G2318,G2177,G1114);
  and AND2_296(G2319,G2185,G816);
  and AND2_297(G2320,G2178,G1115);
  and AND2_298(G2321,G2186,G816);
  and AND2_299(G2322,G2179,G1116);
  and AND2_300(G2323,G2187,G816);
  and AND2_301(G2324,G2180,G1117);
  and AND2_302(G2325,G2188,G816);
  and AND2_303(G2326,G2181,G1118);
  and AND2_304(G2327,G2189,G816);
  and AND2_305(G2328,G2182,G1119);
  and AND2_306(G2329,G2190,G816);
  or OR3_35(G2330,G2198,G2199,G1961);
  or OR3_36(G2331,G2214,G2215,G1977);
  or OR3_37(G2332,G2222,G2223,G1984);
  or OR3_38(G2333,G2230,G2231,G1991);
  or OR3_39(G2334,G2246,G2247,G2007);
  or OR3_40(G2335,G2254,G2255,G2014);
  and AND2_307(G2336,G2256,G1769);
  not NOT_444(G2337,G2263);
  not NOT_445(G2338,G2266);
  not NOT_446(G2339,G2272);
  not NOT_447(G2340,G2269);
  not NOT_448(G2341,G2257);
  not NOT_449(G2342,G2260);
  and AND2_308(G2343,G2313,G1322);
  and AND2_309(G2344,G2311,G1325);
  or OR3_41(G2345,G2314,G2315,G1485);
  or OR2_12(G2346,G2316,G2317);
  or OR2_13(G2347,G2318,G2319);
  or OR2_14(G2348,G2320,G2321);
  or OR2_15(G2349,G2322,G2323);
  or OR2_16(G2350,G2324,G2325);
  or OR2_17(G2351,G2326,G2327);
  or OR2_18(G2352,G2328,G2329);
  and AND2_310(G2353,G2312,G1684);
  or OR2_19(G2354,G2192,G2195);
  nor NOR2_12(G2355,G2192,G2195);
  and AND3_58(G2356,G23,G2200,G1965);
  and AND3_59(G2359,G24,G2200,G1968);
  and AND3_60(G2362,G25,G2204,G1968);
  and AND3_61(G2363,G26,G2204,G1965);
  not NOT_450(G2364,G2204);
  or OR2_20(G2365,G2208,G2211);
  nor NOR2_13(G2368,G2208,G2211);
  or OR2_21(G2369,G2216,G2219);
  nor NOR2_14(G2372,G2216,G2219);
  or OR2_22(G2373,G2224,G2227);
  nor NOR2_15(G2374,G2224,G2227);
  and AND3_62(G2375,G23,G2232,G1995);
  and AND3_63(G2378,G24,G2232,G1998);
  and AND3_64(G2381,G25,G2236,G1998);
  and AND3_65(G2382,G26,G2236,G1995);
  not NOT_451(G2383,G2236);
  or OR2_23(G2384,G2240,G2243);
  nor NOR2_16(G2387,G2240,G2243);
  or OR2_24(G2388,G2248,G2251);
  nor NOR2_17(G2391,G2248,G2251);
  not NOT_452(G2392,G2278);
  and AND2_311(G2393,G1176,G2200);
  not NOT_453(G2396,G2281);
  not NOT_454(G2397,G2284);
  not NOT_455(G2398,G2287);
  not NOT_456(G2399,G2290);
  not NOT_457(G2400,G2296);
  and AND2_312(G2401,G1189,G2232);
  not NOT_458(G2404,G2302);
  not NOT_459(G2405,G2305);
  not NOT_460(G2406,G2308);
  not NOT_461(G2407,G2299);
  not NOT_462(G2408,G2169);
  not NOT_463(G2411,G2169);
  not NOT_464(G2414,G2275);
  not NOT_465(G2415,G2293);
  nand NAND2_84(G2416,G2260,G2341);
  nand NAND2_85(G2417,G2257,G2342);
  nand NAND2_86(G2418,G2266,G2337);
  nand NAND2_87(G2419,G2263,G2338);
  or OR3_42(G2420,G2343,G1473,G1474);
  or OR3_43(G2421,G2344,G1475,G1476);
  and AND2_313(G2422,G2345,G1673);
  and AND2_314(G2423,G2346,G1675);
  and AND2_315(G2424,G2347,G1677);
  and AND2_316(G2425,G2348,G1679);
  and AND2_317(G2426,G2349,G1681);
  and AND2_318(G2427,G2350,G1683);
  and AND2_319(G2428,G2351,G1685);
  and AND2_320(G2429,G2352,G1687);
  and AND2_321(G2430,G2355,G2330);
  or OR3_44(G2436,G2362,G2363,G2364);
  and AND2_322(G2437,G2368,G2331);
  and AND2_323(G2441,G2372,G2332);
  and AND2_324(G2444,G2374,G2333);
  or OR3_45(G2450,G2381,G2382,G2383);
  and AND2_325(G2451,G2387,G2334);
  and AND2_326(G2455,G2391,G2335);
  not NOT_466(G2458,G2354);
  not NOT_467(G2459,G2373);
  nand NAND2_88(G2460,G2416,G2417);
  nand NAND2_89(G2461,G2418,G2419);
  nand NAND2_90(G2462,G2411,G2339);
  not NOT_468(G2463,G2411);
  nand NAND2_91(G2464,G2408,G2340);
  not NOT_469(G2465,G2408);
  and AND2_327(G2466,G2421,G1686);
  and AND2_328(G2467,G2420,G1688);
  or OR2_25(G2468,G2356,G2359);
  nor NOR2_18(G2471,G2356,G2359);
  or OR2_26(G2472,G2375,G2378);
  nor NOR2_19(G2475,G2375,G2378);
  and AND2_329(G2476,G2365,G1184);
  and AND2_330(G2479,G2369,G1184);
  and AND2_331(G2482,G2384,G1193);
  and AND2_332(G2485,G2388,G1193);
  not NOT_470(G2488,G2393);
  not NOT_471(G2491,G2393);
  not NOT_472(G2494,G2401);
  not NOT_473(G2497,G2401);
  nand NAND2_92(G2500,G2272,G2463);
  nand NAND2_93(G2501,G2269,G2465);
  and AND2_333(G2502,G2471,G2436);
  and AND2_334(G2507,G2475,G2450);
  not NOT_474(G2512,G2430);
  not NOT_475(G2515,G2437);
  not NOT_476(G2518,G2441);
  not NOT_477(G2521,G2444);
  not NOT_478(G2524,G2451);
  not NOT_479(G2527,G2455);
  nand NAND2_94(G2530,G2462,G2500);
  nand NAND2_95(G2531,G2464,G2501);
  nand NAND2_96(G2532,G2430,G2468);
  nand NAND2_97(G2533,G2444,G2472);
  not NOT_480(G2534,G2488);
  not NOT_481(G2535,G2491);
  not NOT_482(G2536,G2497);
  not NOT_483(G2537,G2494);
  and AND2_335(G2538,G2468,G1179);
  not NOT_484(G2539,G2479);
  and AND2_336(G2542,G2472,G1184);
  not NOT_485(G2543,G2485);
  not NOT_486(G2546,G2476);
  not NOT_487(G2547,G2485);
  not NOT_488(G2550,G2530);
  not NOT_489(G2551,G2531);
  and AND4_3(G2552,G2430,G2502,G2437,G2441);
  nand NAND3_10(G2556,G2430,G2502,G2365);
  nand NAND4_1(G2557,G2369,G2502,G2437,G2430);
  and AND4_4(G2558,G2444,G2507,G2451,G2455);
  nand NAND3_11(G2561,G2444,G2507,G2384);
  nand NAND4_2(G2562,G2388,G2507,G2451,G2444);
  not NOT_490(G2563,G2502);
  not NOT_491(G2566,G2507);
  not NOT_492(G2569,G2538);
  not NOT_493(G2570,G2542);
  not NOT_494(G2571,G2512);
  not NOT_495(G2574,G2512);
  not NOT_496(G2577,G2515);
  not NOT_497(G2580,G2515);
  not NOT_498(G2583,G2518);
  not NOT_499(G2586,G2518);
  not NOT_500(G2589,G2521);
  not NOT_501(G2592,G2521);
  not NOT_502(G2595,G2524);
  not NOT_503(G2598,G2524);
  not NOT_504(G2601,G2527);
  not NOT_505(G2604,G2527);
  nand NAND4_3(G2607,G2458,G2532,G2556,G2557);
  nand NAND4_4(G2610,G2459,G2533,G2561,G2562);
  not NOT_506(G2613,G2547);
  nand NAND2_98(G2614,G2574,G2392);
  nand NAND2_99(G2615,G2580,G2397);
  nand NAND2_100(G2616,G2586,G2399);
  nand NAND2_101(G2617,G2592,G2400);
  nand NAND2_102(G2618,G2598,G2404);
  nand NAND2_103(G2619,G2604,G2406);
  not NOT_507(G2620,G2552);
  not NOT_508(G2623,G2574);
  not NOT_509(G2624,G2577);
  nand NAND2_104(G2625,G2577,G2396);
  not NOT_510(G2626,G2580);
  not NOT_511(G2627,G2583);
  nand NAND2_105(G2628,G2583,G2398);
  not NOT_512(G2629,G2586);
  not NOT_513(G2630,G2592);
  not NOT_514(G2631,G2598);
  not NOT_515(G2632,G2601);
  nand NAND2_106(G2633,G2601,G2405);
  not NOT_516(G2634,G2604);
  not NOT_517(G2635,G2595);
  nand NAND2_107(G2636,G2595,G2407);
  and AND2_337(G2637,G2558,G1433);
  not NOT_518(G2638,G2571);
  nand NAND2_108(G2639,G2571,G2414);
  not NOT_519(G2640,G2563);
  not NOT_520(G2643,G2563);
  not NOT_521(G2646,G2589);
  nand NAND2_109(G2647,G2589,G2415);
  not NOT_522(G2648,G2566);
  not NOT_523(G2651,G2566);
  nand NAND2_110(G2654,G2552,G2610);
  not NOT_524(G2655,G2607);
  nand NAND2_111(G2656,G2278,G2623);
  nand NAND2_112(G2657,G2284,G2626);
  nand NAND2_113(G2658,G2290,G2629);
  nand NAND2_114(G2659,G2296,G2630);
  nand NAND2_115(G2660,G2302,G2631);
  nand NAND2_116(G2661,G2308,G2634);
  nand NAND2_117(G2662,G2281,G2624);
  nand NAND2_118(G2663,G2287,G2627);
  nand NAND2_119(G2664,G2305,G2632);
  nand NAND2_120(G2665,G2299,G2635);
  and AND2_338(G2666,G2610,G1193);
  or OR2_27(G2669,G2336,G2637);
  nand NAND2_121(G2673,G2275,G2638);
  nand NAND2_122(G2674,G2293,G2646);
  and AND2_339(G2675,G2654,G2655);
  nand NAND2_123(G2676,G2656,G2614);
  nand NAND2_124(G2677,G2643,G2535);
  nand NAND2_125(G2678,G2657,G2615);
  nand NAND2_126(G2679,G2658,G2616);
  nand NAND2_127(G2680,G2659,G2617);
  nand NAND2_128(G2681,G2651,G2536);
  nand NAND2_129(G2682,G2660,G2618);
  nand NAND2_130(G2683,G2661,G2619);
  not NOT_525(G2684,G2640);
  nand NAND2_131(G2685,G2640,G2534);
  not NOT_526(G2686,G2643);
  nand NAND2_132(G2687,G2662,G2625);
  nand NAND2_133(G2690,G2663,G2628);
  not NOT_527(G2693,G2651);
  nand NAND2_134(G2694,G2664,G2633);
  not NOT_528(G2697,G2648);
  nand NAND2_135(G2698,G2648,G2537);
  nand NAND2_136(G2699,G2665,G2636);
  nand NAND2_137(G2705,G2673,G2639);
  nand NAND2_138(G2708,G2674,G2647);
  not NOT_529(G2711,G2676);
  nand NAND2_139(G2712,G2491,G2686);
  not NOT_530(G2713,G2678);
  not NOT_531(G2714,G2679);
  not NOT_532(G2715,G2680);
  nand NAND2_140(G2716,G2497,G2693);
  not NOT_533(G2717,G2682);
  not NOT_534(G2718,G2683);
  nand NAND2_141(G2719,G2488,G2684);
  nand NAND2_142(G2720,G2494,G2697);
  not NOT_535(G2721,G2666);
  not NOT_536(G2728,G2669);
  not NOT_537(G2733,G2666);
  and AND2_340(G2736,G47,G2669);
  and AND2_341(G2739,G2711,G1399);
  nand NAND2_143(G2740,G2712,G2677);
  and AND2_342(G2741,G2713,G1401);
  and AND2_343(G2742,G2714,G1402);
  and AND2_344(G2743,G2715,G1403);
  nand NAND2_144(G2744,G2716,G2681);
  and AND2_345(G2745,G2717,G1405);
  and AND2_346(G2746,G2718,G1406);
  nand NAND2_145(G2747,G2719,G2685);
  not NOT_538(G2750,G2687);
  not NOT_539(G2753,G2687);
  not NOT_540(G2759,G2690);
  not NOT_541(G2763,G2690);
  nand NAND2_146(G2768,G2720,G2698);
  not NOT_542(G2773,G2694);
  and AND2_347(G2778,G2699,G2543);
  not NOT_543(G2779,G2705);
  not NOT_544(G2780,G2708);
  and AND2_348(G2781,G47,G2694);
  not NOT_545(G2784,G2699);
  nor NOR3_9(G2787,G2422,G2739,G1807);
  not NOT_546(G2788,G2740);
  nor NOR3_10(G2789,G2424,G2741,G1809);
  nor NOR3_11(G2790,G2425,G2742,G1810);
  nor NOR3_12(G2791,G2426,G2743,G2191);
  not NOT_547(G2792,G2744);
  nor NOR3_13(G2793,G2428,G2745,G2466);
  nor NOR3_14(G2794,G2429,G2746,G2467);
  and AND2_349(G2795,G2721,G2620);
  and AND2_350(G2796,G2728,G2620);
  or OR2_28(G2799,G2482,G2778);
  not NOT_548(G2803,G2736);
  not NOT_549(G2804,G2721);
  not NOT_550(G2805,G2721);
  not NOT_551(G2808,G2733);
  and AND2_351(G2809,G2788,G1400);
  and AND2_352(G2810,G2792,G1404);
  not NOT_552(G2811,G2747);
  or OR2_29(G2816,G2607,G2795);
  and AND3_66(G2820,G2728,G2763,G2753);
  and AND2_353(G2821,G2728,G2759);
  and AND3_67(G2822,G2773,G2699,G2768);
  and AND2_354(G2823,G2773,G2699);
  and AND2_355(G2826,G2721,G2759);
  nand NAND2_147(G2827,G2753,G2539);
  nand NAND3_12(G2828,G2753,G2763,G2721);
  nand NAND2_148(G2829,G2768,G2482);
  nand NAND3_13(G2830,G2768,G2699,G2543);
  nand NAND2_149(G2831,G2784,G2613);
  not NOT_553(G2832,G2784);
  and AND3_68(G2833,G47,G2669,G2804);
  and AND2_356(G2836,G2787,G1771);
  and AND2_357(G2839,G2789,G1775);
  and AND2_358(G2842,G2790,G1777);
  and AND2_359(G2845,G2791,G1779);
  and AND2_360(G2848,G2793,G1783);
  and AND2_361(G2851,G2794,G1785);
  not NOT_554(G2854,G2747);
  not NOT_555(G2857,G2753);
  not NOT_556(G2860,G2759);
  not NOT_557(G2863,G2768);
  not NOT_558(G2866,G2781);
  not NOT_559(G2869,G2781);
  and AND2_362(G2872,G2773,G2773);
  nor NOR3_15(G2875,G2423,G2809,G1808);
  nor NOR3_16(G2876,G2427,G2810,G2353);
  and AND2_363(G2877,G47,G2821);
  and AND2_364(G2880,G47,G2822);
  nand NAND2_150(G2883,G2547,G2832);
  not NOT_560(G2884,G2799);
  not NOT_561(G2887,G2796);
  nand NAND3_14(G2890,G2546,G2827,G2828);
  or OR2_30(G2893,G2479,G2826);
  nand NAND3_15(G2896,G2570,G2829,G2830);
  not NOT_562(G2899,G2799);
  and AND2_365(G2902,G47,G2820);
  or OR2_31(G2905,G2833,G2805);
  and AND4_5(G2906,G2728,G2811,G2753,G2763);
  nand NAND2_151(G2909,G2811,G2476);
  nand NAND3_16(G2910,G2811,G2750,G2539);
  nand NAND4_5(G2911,G2811,G2750,G2763,G2721);
  not NOT_563(G2912,G2857);
  nand NAND2_152(G2913,G2831,G2883);
  not NOT_564(G2916,G2866);
  not NOT_565(G2917,G2869);
  nand NAND2_153(G2918,G2872,G883);
  not NOT_566(G2919,G2872);
  not NOT_567(G2920,G2816);
  nor NOR2_20(G2923,G2833,G2805);
  and AND2_366(G2926,G2875,G1773);
  and AND2_367(G2929,G2876,G1781);
  not NOT_568(G2932,G2816);
  not NOT_569(G2935,G2854);
  not NOT_570(G2936,G2860);
  nand NAND2_154(G2937,G2860,G2808);
  not NOT_571(G2938,G2863);
  and AND2_368(G2939,G47,G2823);
  not NOT_572(G2942,G2884);
  and AND2_369(G2943,G2799,G2884);
  and AND2_370(G2944,G2905,G1056);
  nand NAND4_6(G2947,G2569,G2909,G2910,G2911);
  not NOT_573(G2950,G2887);
  not NOT_574(G2951,G2902);
  not NOT_575(G2952,G2893);
  nand NAND2_155(G2953,G2893,G2912);
  not NOT_576(G2954,G2896);
  nand NAND2_156(G2955,G2896,G2780);
  nand NAND2_157(G2956,G663,G2919);
  not NOT_577(G2957,G2890);
  nand NAND2_158(G2958,G2890,G2935);
  nand NAND2_159(G2959,G2733,G2936);
  not NOT_578(G2960,G2899);
  nand NAND2_160(G2961,G2899,G2938);
  not NOT_579(G2962,G2877);
  not NOT_580(G2965,G2877);
  not NOT_581(G2968,G2880);
  not NOT_582(G2971,G2880);
  and AND3_69(G2974,G47,G2823,G2942);
  and AND2_371(G2975,G47,G2906);
  nand NAND2_161(G2978,G2857,G2952);
  nand NAND2_162(G2979,G2708,G2954);
  not NOT_583(G2980,G2939);
  nand NAND2_163(G2981,G2918,G2956);
  not NOT_584(G2984,G2920);
  and AND2_372(G2985,G2816,G2920);
  not NOT_585(G2986,G2923);
  not NOT_586(G2990,G2932);
  not NOT_587(G2991,G2906);
  nand NAND2_164(G2994,G2854,G2957);
  nand NAND2_165(G2995,G2863,G2960);
  nand NAND2_166(G2996,G2937,G2959);
  not NOT_588(G2999,G2913);
  not NOT_589(G3002,G2913);
  or OR3_46(G3005,G1796,G2944,G1799);
  nor NOR3_17(G3006,G1796,G2944,G1799);
  nand NAND2_167(G3007,G2978,G2953);
  not NOT_590(G3010,G2962);
  not NOT_591(G3011,G2965);
  nand NAND2_168(G3012,G2979,G2955);
  not NOT_592(G3015,G2968);
  not NOT_593(G3016,G2971);
  and AND3_70(G3017,G47,G2796,G2984);
  not NOT_594(G3018,G2947);
  not NOT_595(G3021,G2947);
  nand NAND2_169(G3024,G2994,G2958);
  nand NAND2_170(G3027,G2995,G2961);
  not NOT_596(G3030,G3006);
  nand NAND2_171(G3031,G2991,G2950);
  not NOT_597(G3032,G2991);
  not NOT_598(G3033,G2996);
  nand NAND2_172(G3034,G2996,G2803);
  not NOT_599(G3035,G2999);
  nand NAND2_173(G3036,G2999,G2916);
  not NOT_600(G3037,G3002);
  nand NAND2_174(G3038,G3002,G2917);
  nor NOR2_21(G3039,G3017,G2985);
  and AND2_373(G3042,G2981,G1303);
  and AND2_374(G3045,G2981,G1784);
  not NOT_601(G3048,G2975);
  not NOT_602(G3051,G2975);
  not NOT_603(G3054,G2986);
  nand NAND2_175(G3057,G2887,G3032);
  not NOT_604(G3058,G3021);
  nand NAND2_176(G3059,G3021,G2779);
  not NOT_605(G3060,G3024);
  nand NAND2_177(G3061,G3024,G2951);
  nand NAND2_178(G3062,G2736,G3033);
  not NOT_606(G3063,G3027);
  nand NAND2_179(G3064,G3027,G2980);
  nand NAND2_180(G3065,G2866,G3035);
  nand NAND2_181(G3066,G2869,G3037);
  not NOT_607(G3067,G3018);
  nand NAND2_182(G3068,G3018,G2990);
  not NOT_608(G3069,G3007);
  not NOT_609(G3072,G3007);
  not NOT_610(G3075,G3012);
  not NOT_611(G3078,G3012);
  nand NAND2_183(G3081,G3031,G3057);
  nand NAND2_184(G3082,G2705,G3058);
  not NOT_612(G3083,G3048);
  not NOT_613(G3084,G3051);
  nand NAND2_185(G3085,G2902,G3060);
  nand NAND2_186(G3086,G3062,G3034);
  nand NAND2_187(G3089,G2939,G3063);
  nand NAND2_188(G3090,G3065,G3036);
  nand NAND2_189(G3094,G3066,G3038);
  not NOT_614(G3095,G3039);
  not NOT_615(G3099,G3054);
  or OR3_47(G3100,G3042,G3045,G2851);
  nor NOR3_18(G3103,G3042,G3045,G2851);
  nand NAND2_190(G3106,G2932,G3067);
  nand NAND2_191(G3107,G3082,G3059);
  nand NAND2_192(G3110,G3085,G3061);
  not NOT_616(G3114,G3069);
  nand NAND2_193(G3115,G3069,G3010);
  not NOT_617(G3116,G3072);
  nand NAND2_194(G3117,G3072,G3011);
  not NOT_618(G3118,G3075);
  nand NAND2_195(G3119,G3075,G3015);
  not NOT_619(G3120,G3078);
  nand NAND2_196(G3121,G3078,G3016);
  nand NAND2_197(G3122,G3089,G3064);
  nand NAND2_198(G3126,G3106,G3068);
  and AND2_375(G3129,G47,G3081);
  not NOT_620(G3132,G3094);
  not NOT_621(G3135,G3103);
  nand NAND2_199(G3136,G2962,G3114);
  nand NAND2_200(G3137,G2965,G3116);
  nand NAND2_201(G3138,G2968,G3118);
  nand NAND2_202(G3139,G2971,G3120);
  and AND2_376(G3140,G3086,G1299);
  and AND2_377(G3143,G3086,G1776);
  and AND2_378(G3146,G3090,G1302);
  not NOT_622(G3149,G3095);
  and AND2_379(G3152,G3090,G2923);
  not NOT_623(G3155,G3100);
  not NOT_624(G3158,G3126);
  not NOT_625(G3159,G3129);
  nand NAND2_203(G3160,G3136,G3115);
  nand NAND2_204(G3164,G3137,G3117);
  nand NAND2_205(G3165,G3138,G3119);
  nand NAND2_206(G3168,G3139,G3121);
  nand NAND2_207(G3169,G3132,G3099);
  not NOT_626(G3170,G3132);
  and AND2_380(G3171,G3110,G1297);
  and AND2_381(G3174,G3122,G1301);
  not NOT_627(G3177,G3107);
  not NOT_628(G3180,G3107);
  not NOT_629(G3183,G3110);
  not NOT_630(G3186,G3122);
  nand NAND2_208(G3189,G3129,G3158);
  nand NAND2_209(G3190,G3126,G3159);
  not NOT_631(G3191,G3168);
  not NOT_632(G3192,G3149);
  not NOT_633(G3193,G3152);
  nand NAND2_210(G3194,G3054,G3170);
  or OR3_48(G3195,G3140,G3143,G2842);
  nor NOR3_19(G3199,G3140,G3143,G2842);
  not NOT_634(G3202,G3155);
  not NOT_635(G3203,G3164);
  nand NAND2_211(G3206,G3189,G3190);
  not NOT_636(G3207,G3177);
  nand NAND2_212(G3208,G3177,G3083);
  not NOT_637(G3209,G3180);
  nand NAND2_213(G3210,G3180,G3084);
  nor NOR2_22(G3211,G3191,G2986);
  and AND4_6(G3212,G3090,G3122,G3165,G2986);
  not NOT_638(G3213,G3183);
  not NOT_639(G3214,G3186);
  nand NAND2_214(G3215,G3186,G3193);
  nand NAND2_215(G3216,G3194,G3169);
  and AND2_382(G3217,G3160,G1298);
  and AND2_383(G3220,G3165,G1300);
  and AND2_384(G3223,G3160,G3039);
  not NOT_640(G3226,G3199);
  and AND2_385(G3227,G3206,G1353);
  nand NAND2_216(G3230,G3048,G3207);
  nand NAND2_217(G3231,G3051,G3209);
  or OR2_32(G3232,G3211,G3212);
  nand NAND2_218(G3233,G3203,G3192);
  not NOT_641(G3234,G3203);
  nand NAND2_219(G3235,G3152,G3214);
  not NOT_642(G3236,G3216);
  not NOT_643(G3237,G3195);
  not NOT_644(G3240,G3195);
  nand NAND2_220(G3243,G3230,G3208);
  nand NAND2_221(G3246,G3231,G3210);
  nand NAND2_222(G3247,G3223,G3213);
  not NOT_645(G3248,G3223);
  nand NAND2_223(G3249,G3149,G3234);
  nand NAND2_224(G3250,G3235,G3215);
  and AND2_386(G3251,G3232,G1778);
  and AND2_387(G3254,G3236,G1782);
  or OR3_49(G3257,G1802,G1524,G3227);
  nor NOR3_20(G3258,G1802,G1524,G3227);
  not NOT_646(G3259,G3246);
  nand NAND2_225(G3260,G3183,G3248);
  nand NAND2_226(G3261,G3249,G3233);
  and AND2_388(G3262,G3250,G1780);
  not NOT_647(G3265,G3237);
  not NOT_648(G3266,G3240);
  not NOT_649(G3267,G3258);
  nor NOR2_23(G3268,G3259,G3095);
  and AND4_7(G3269,G3160,G3110,G3243,G3095);
  nand NAND2_227(G3270,G3247,G3260);
  not NOT_650(G3271,G3261);
  and AND2_389(G3272,G3243,G1296);
  or OR3_50(G3275,G3220,G3251,G2845);
  nor NOR3_21(G3278,G3220,G3251,G2845);
  or OR3_51(G3281,G3146,G3254,G2848);
  nor NOR3_22(G3284,G3146,G3254,G2848);
  or OR2_33(G3287,G3268,G3269);
  and AND2_390(G3288,G3270,G1772);
  and AND2_391(G3291,G3271,G1774);
  or OR3_52(G3294,G3174,G3262,G2929);
  nor NOR3_23(G3297,G3174,G3262,G2929);
  not NOT_651(G3300,G3278);
  not NOT_652(G3301,G3284);
  and AND2_392(G3302,G3287,G1770);
  not NOT_653(G3305,G3281);
  not NOT_654(G3308,G3275);
  not NOT_655(G3311,G3297);
  or OR3_53(G3312,G3171,G3288,G2926);
  nor NOR3_24(G3317,G3171,G3288,G2926);
  or OR3_54(G3320,G3217,G3291,G2839);
  nor NOR3_25(G3323,G3217,G3291,G2839);
  and AND4_8(G3326,G3103,G3284,G3297,G3278);
  not NOT_656(G3329,G3294);
  or OR3_55(G3332,G3272,G3302,G2836);
  nor NOR3_26(G3337,G3272,G3302,G2836);
  nand NAND2_228(G3340,G3305,G3202);
  not NOT_657(G3341,G3305);
  not NOT_658(G3342,G3308);
  not NOT_659(G3343,G3323);
  nand NAND2_229(G3344,G3155,G3341);
  not NOT_660(G3345,G3329);
  nand NAND2_230(G3346,G3329,G3342);
  not NOT_661(G3347,G3320);
  and AND2_393(G3350,G3312,G884);
  not NOT_662(G3353,G3312);
  nand NAND2_231(G3356,G3340,G3344);
  nand NAND2_232(G3359,G3308,G3345);
  and AND2_394(G3360,G884,G3332);
  and AND4_9(G3363,G3199,G3323,G3317,G3337);
  and AND3_71(G3366,G3317,G3337,G887);
  not NOT_663(G3367,G3332);
  nand NAND2_233(G3370,G3359,G3346);
  not NOT_664(G3373,G3347);
  not NOT_665(G3376,G3347);
  not NOT_666(G3379,G3353);
  not NOT_667(G3380,G3350);
  not NOT_668(G3383,G3350);
  and AND2_395(G3386,G3326,G3363);
  and AND2_396(G3387,G3326,G3363);
  not NOT_669(G3388,G3356);
  not NOT_670(G3391,G3356);
  not NOT_671(G3394,G3367);
  nand NAND2_234(G3395,G3367,G3379);
  not NOT_672(G3396,G3360);
  not NOT_673(G3399,G3360);
  nor NOR2_24(G3402,G3366,G3387);
  nand NAND2_235(G3403,G3373,G3265);
  not NOT_674(G3404,G3373);
  nand NAND2_236(G3405,G3376,G3266);
  not NOT_675(G3406,G3376);
  not NOT_676(G3407,G3380);
  not NOT_677(G3408,G3383);
  not NOT_678(G3409,G3370);
  not NOT_679(G3412,G3370);
  nand NAND2_237(G3415,G3353,G3394);
  and AND2_397(G3416,G27,G3402);
  not NOT_680(G3417,G3388);
  not NOT_681(G3418,G3391);
  nand NAND2_238(G3419,G3237,G3404);
  nand NAND2_239(G3420,G3240,G3406);
  not NOT_682(G3421,G3396);
  nand NAND2_240(G3422,G3396,G3407);
  nand NAND2_241(G3423,G3399,G3408);
  not NOT_683(G3424,G3399);
  nand NAND2_242(G3425,G3395,G3415);
  nand NAND2_243(G3428,G3409,G3417);
  not NOT_684(G3429,G3409);
  nand NAND2_244(G3430,G3412,G3418);
  not NOT_685(G3431,G3412);
  nand NAND2_245(G3432,G3403,G3419);
  nand NAND2_246(G3436,G3405,G3420);
  nand NAND2_247(G3437,G3380,G3421);
  nand NAND2_248(G3438,G3383,G3424);
  nand NAND2_249(G3439,G3388,G3429);
  nand NAND2_250(G3440,G3391,G3431);
  not NOT_686(G3441,G3436);
  not NOT_687(G3444,G3425);
  nand NAND2_251(G3445,G3437,G3422);
  nand NAND2_252(G3448,G3438,G3423);
  nand NAND2_253(G3449,G3428,G3439);
  nand NAND2_254(G3452,G3430,G3440);
  not NOT_688(G3453,G3448);
  not NOT_689(G3456,G3432);
  and AND3_72(G3459,G3432,G3445,G1436);
  and AND3_73(G3460,G3441,G3445,G1439);
  not NOT_690(G3461,G3452);
  not NOT_691(G3464,G3456);
  nand NAND2_255(G3465,G3456,G3444);
  and AND3_74(G3466,G3432,G3453,G1439);
  and AND3_75(G3467,G3441,G3453,G1436);
  not NOT_692(G3468,G3449);
  not NOT_693(G3471,G3449);
  nand NAND2_256(G3474,G3425,G3464);
  or OR4_0(G3475,G3459,G3466,G3460,G3467);
  not NOT_694(G3478,G3461);
  not NOT_695(G3481,G3461);
  nand NAND2_257(G3484,G3474,G3465);
  not NOT_696(G3487,G3471);
  not NOT_697(G3488,G3468);
  not NOT_698(G3489,G3481);
  not NOT_699(G3490,G3478);
  not NOT_700(G3491,G3475);
  not NOT_701(G3494,G3475);
  not NOT_702(G3497,G3484);
  not NOT_703(G3500,G3484);
  nand NAND2_258(G3503,G3491,G3490);
  nand NAND2_259(G3504,G3494,G3489);
  not NOT_704(G3505,G3494);
  not NOT_705(G3506,G3491);
  nand NAND2_260(G3507,G3497,G3488);
  nand NAND2_261(G3508,G3500,G3487);
  nand NAND2_262(G3509,G3478,G3506);
  nand NAND2_263(G3510,G3481,G3505);
  not NOT_706(G3511,G3500);
  not NOT_707(G3512,G3497);
  nand NAND2_264(G3513,G3468,G3512);
  nand NAND2_265(G3514,G3471,G3511);
  nand NAND2_266(G3515,G3509,G3503);
  nand NAND2_267(G3516,G3510,G3504);
  nand NAND2_268(G3517,G3507,G3513);
  nand NAND2_269(G3518,G3508,G3514);
  not NOT_708(G3519,G928);
  not NOT_709(G3520,G1004);
  nand NAND2_270(G3521,G1786,G1811);
  nand NAND2_271(G3522,G2460,G2461);
  nand NAND2_272(G3523,G2550,G2551);
  and AND2_398(G3524,G2558,G2552);
  not NOT_710(G3525,G2675);
  or OR2_34(G3526,G2974,G2943);
  and AND2_399(G3527,G3005,G3030);
  and AND2_400(G3528,G3100,G3135);
  and AND2_401(G3529,G3195,G3226);
  and AND2_402(G3530,G3257,G3267);
  and AND2_403(G3531,G3275,G3300);
  and AND2_404(G3532,G3281,G3301);
  and AND2_405(G3533,G3294,G3311);
  and AND2_406(G3534,G3312,G3312);
  and AND2_407(G3535,G3332,G3332);
  and AND2_408(G3536,G3320,G3343);
  not NOT_711(G3537,G3386);
  not NOT_712(G3538,G3416);
  and AND2_409(G3539,G3515,G3516);
  nand NAND2_273(G3540,G3517,G3518);

endmodule
